// Verilog netlist created by TD v4.4.433
// Mon May 13 08:51:04 2019

`timescale 1ns / 1ps
module ImgROM  // al_ip/ROM.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [14:0] addra;  // al_ip/ROM.v(18)
  input clka;  // al_ip/ROM.v(19)
  input rsta;  // al_ip/ROM.v(20)
  output [7:0] doa;  // al_ip/ROM.v(16)

  wire [0:1] addra_piped;
  wire  \inst_doa_mux_b0/B0_0 ;
  wire  \inst_doa_mux_b0/B0_1 ;
  wire  \inst_doa_mux_b1/B0_0 ;
  wire  \inst_doa_mux_b1/B0_1 ;
  wire  \inst_doa_mux_b2/B0_0 ;
  wire  \inst_doa_mux_b2/B0_1 ;
  wire  \inst_doa_mux_b3/B0_0 ;
  wire  \inst_doa_mux_b3/B0_1 ;
  wire  \inst_doa_mux_b4/B0_0 ;
  wire  \inst_doa_mux_b4/B0_1 ;
  wire  \inst_doa_mux_b5/B0_0 ;
  wire  \inst_doa_mux_b5/B0_1 ;
  wire  \inst_doa_mux_b6/B0_0 ;
  wire  \inst_doa_mux_b6/B0_1 ;
  wire  \inst_doa_mux_b7/B0_0 ;
  wire  \inst_doa_mux_b7/B0_1 ;
  wire inst_doa_i0_000;
  wire inst_doa_i0_001;
  wire inst_doa_i0_002;
  wire inst_doa_i0_003;
  wire inst_doa_i0_004;
  wire inst_doa_i0_005;
  wire inst_doa_i0_006;
  wire inst_doa_i0_007;
  wire inst_doa_i1_000;
  wire inst_doa_i1_001;
  wire inst_doa_i1_002;
  wire inst_doa_i1_003;
  wire inst_doa_i1_004;
  wire inst_doa_i1_005;
  wire inst_doa_i1_006;
  wire inst_doa_i1_007;
  wire inst_doa_i2_000;
  wire inst_doa_i2_001;
  wire inst_doa_i2_002;
  wire inst_doa_i2_003;
  wire inst_doa_i2_004;
  wire inst_doa_i2_005;
  wire inst_doa_i2_006;
  wire inst_doa_i2_007;
  wire inst_doa_i3_000;
  wire inst_doa_i3_001;
  wire inst_doa_i3_002;
  wire inst_doa_i3_003;
  wire inst_doa_i3_004;
  wire inst_doa_i3_005;
  wire inst_doa_i3_006;
  wire inst_doa_i3_007;

  reg_sr_as_w1 addra_pipe_b0 (
    .clk(clka),
    .d(addra[13]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[0]));
  reg_sr_as_w1 addra_pipe_b1 (
    .clk(clka),
    .d(addra[14]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[1]));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFCEA9AF7E9AAAAAAAAACBBFC2AE75BEEFBBFCFAAAAAAAAAAAAAAAAAAAEBD039),
    .INIT_01(256'hFFABFBAD360FFFFFFFFFBF8B52FFB3FE2EB8FEEFFFFFFFFAFEFFEFFFF9CD1F7D),
    .INIT_02(256'hFF8FBEBEEEAFFFFFFFFEBF8A3AE24D2E6AA2ABAFFFFEBBB9E0EAAD783F9F3F82),
    .INIT_03(256'hFF9FAFA7BDAFFFFFFFFFDF9C0AE9E2AE6A9EDFFAFFFAF37B9750725982FEBB1F),
    .INIT_04(256'hFF8EDAF6C8BFFFFFFFFF0B8DEA8BEF4E22CEFFFAFFE83986BF3FEDAFABEE90FB),
    .INIT_05(256'hFF8E2FFC8AEFFFFFEAF92B8C6ED181DEE36E7FFFFFE75BFE083383AFEFFB27FF),
    .INIT_06(256'hFF9E6AEEDBBFFFFFEAFEFEB5AE3BFA9AE6A9FFFFFFEEFE3576ED3AFFFEEA7FFF),
    .INIT_07(256'hFF8FB2FD7BFFFFFFEAFFBA76BAACB456A1AEBFFFFFFBBA73AF4EBFFFFE90EFFF),
    .INIT_08(256'hFFABFFFF6FFFEAFFEAAC2F21A83BFC13A3E6FFFFBAE6E6EFA5ABFFFFFFBBF924),
    .INIT_09(256'hFFEBE3FF8FFFFEBFEAA4FE17A58D3D85BFF7FFFFFDFCBFAC2ABFEBFFFFAE95C3),
    .INIT_0A(256'hFFCADEEE9BFFFCAFEAF2FE4ABE4EEE3EFFDBFFFA932AEB0EBFFAABFFFEBBC001),
    .INIT_0B(256'hFF92A7EEEFFFE86BEBFFFE268DFE5F29BFBBFBFBAEFBB5AFFFFEABFEBFE505AA),
    .INIT_0C(256'hFFE784ADAFFFCAE6BFF9BEA7692FFBB33E2BFAE8BFFD7EAAAAAABFFFFFEDBFFF),
    .INIT_0D(256'hFFEBA6EEFEBF8DFDAFBDBA0E7E5AEF8D3E6BFA8EFFED40000153AAFFFFFBFFFF),
    .INIT_0E(256'hFFCABCEFA6EBE72E9EAFAA6EF6E416D33CBAE9ABFFFAAAAAAAAEC5AAAFFEFFFF),
    .INIT_0F(256'hFFE3BEB8BB2BE8A2F6DFA9DC90FFFAD4F9AFB6BFFFFEFFFFFFFFAAE4ABFBA4FF),
    .INIT_10(256'hCECEE4B9BE86AAEABF73A9F8F8251151E6AB7FFC2AFFFFFFFFFFFFAAC6AAED4F),
    .INIT_11(256'hEAB0A8E8BFE96A6BFABFB97EE8FC1FD0E2AEB0A30CBFFFFFFFFFFFFFFB5ABBA7),
    .INIT_12(256'h7DADEE29BFFFC6DEBC66BB32D0C3A2B3AA877272A6EF056FFFFFFFFFFAF86ADA),
    .INIT_13(256'h5F1DBBCAFFFFFB13260ABEB209B59125CAA91F13C1A901CBB06FFFFFF0107AE8),
    .INIT_14(256'h9696EDBF6FFFFFBF8E3AFC7F334E9744B66C645B19DD707FCAD96AAABAAAAAFA),
    .INIT_15(256'hC7E8BEB76FFFEFEFE6FFA95D1E24529E3F38EE9ABAEF907FF8505F3ABFFEBFFA),
    .INIT_16(256'hF3EC7B5EBBFFFEBCAF3FADAE4BFFEFF17BAEBFFEABEF3943FFFFB1CF5BBFFFFF),
    .INIT_17(256'hFB6E6BDDCBFFFFCC1B3FAEBDAFFFFFFEAFEEFFFFFFEAE1823FFFFFA50A2EAFFF),
    .INIT_18(256'hFFAAAE0E8BFFFCB11BDFAA312FFFFFFEAAAEFFFFFFFABB8EE3FFFFEAE81CFAFB),
    .INIT_19(256'hFFAEFA8A6BFFFB3DF89F8E2DAEBFFFFEAABFFFFFFFFFFC4F8FFFFFFFFFF3B3AA),
    .INIT_1A(256'hFF5FFEAEEBFFE5CAE8BF5AE2AEBFFFFFFABFFFFFFFFEBE5A30FFFFFFFFFEADCA),
    .INIT_1B(256'hFFE6FFEE86FFE23ABEDA08C8AEFFFFFFFEBFFFFEAFEABA6C1BFFFFFFFFFFECE1),
    .INIT_1C(256'hFFE1ABE2E6FF3F6FFE4A5CA3FFFFFFFFFFFFFFFFAEEAA8C68CFFFFFFFFFFFFBE),
    .INIT_1D(256'hFFF2BFE6FFFE2DFFFFFADDBAAFFFFFFFFFFFFFFFFEFAAE3AB06FFFFFFFFFFFFB),
    .INIT_1E(256'hE7F92FE2FBFDE4EFFEBB9B9ABFFFFFFFFFFFFFFFFB62A61E792FFFFFFFFFFFFF),
    .INIT_1F(256'h9B2DFEA7FBFE7B6FFCA9D75EFFFFFFFFFFFFFFFFEBA8A057998BFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_000000_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n63,addra[14:13]}),
    .dia({open_n67,open_n68,open_n69,open_n70,open_n71,open_n72,open_n73,1'b0,open_n74}),
    .rsta(rsta),
    .doa({open_n89,open_n90,open_n91,open_n92,open_n93,open_n94,open_n95,open_n96,inst_doa_i0_000}));
  // address_offset=0;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFBEABBC742AAAAAAAAA92B50AAF5ABED6BB542AAAAAAAAAAAAAAAAAAABEEAEE),
    .INIT_01(256'hFFBBFA0F6B7FFFFFFFFFBFB51EF856BED6BA58AFFFFFFFFAABAAAAAAAA0EAFEE),
    .INIT_02(256'hFF8BBEBB6BEFFFFFFFFE7BB51AED66AE92AD22AFFFFEBAEA44FAA9112F95FB63),
    .INIT_03(256'hFF8BAF9738BFFFFFFFFEDBA47AFB1AFE92B48BFAFFFAAC2AC4EF82AC2EAAAAEF),
    .INIT_04(256'hFF9AFAE67A2FFFFFFFFEEBA42AA535BE9AE6AFFAFFEB692EFE9EBC6AABEEFDFF),
    .INIT_05(256'hFF9ACBE53AEFFFFFEAFAEBA0AEBE12CA5A96FFFFFFEB6AAA9AA46FAFEFFA6FFF),
    .INIT_06(256'hFF8AFAEBABBFFFFFEAF8EE95AE9C5D7A5A57BFFFFFEEAAC7B446FAFFFEEB3FFF),
    .INIT_07(256'hFF8BBEFB1BFFFFFFEAFA2AD1BAF015AE5E56BFFFFFFA8E7405FEBFFFFEA8BFFF),
    .INIT_08(256'hFFBBB6FE8BFFEAFFEAAEEFD2AAC314B2595AFFFFBAA8A1454BABFFFFFF9AED4F),
    .INIT_09(256'hFFABB6FE5BFFFEBFEAAFBED3A9A5150B555FFFFFEA7D5556EABFEBFFFFAABB13),
    .INIT_0A(256'hFFBA8BEEABFFFFAFEAE7BE82B7259540556BFFFAB35055BEBFFAABFFFEBAFFFE),
    .INIT_0B(256'hFFEE9AEEEFFFEAEBEBEDBEBEA6941554157BFBFA30515BAFFFFEABFEBFEA11FF),
    .INIT_0C(256'hFFEEBFAEAFFFFA5EBFEFBE7ED375310E95ABFAEB5556EAAAAAAABFFFFFEF7FFF),
    .INIT_0D(256'hFFE2A9AD7ABFB792AFAABA4A9E98714E95EBFAB55556AAAAAAAFAAFFFFFB9FFF),
    .INIT_0E(256'hBFCFA9AD5AABE8E53AABAA4A5D41805596BAEB155555555555516BAAAFFEE7FF),
    .INIT_0F(256'h9FCEA6FA55EBEA4C5AAAABBB5A574C5657AFBD55555555555555554BABFBA4FF),
    .INIT_10(256'h8FF6EBBA556EAA5015C6AABA6F592C925EAB955685555555555555556EAAE8FF),
    .INIT_11(256'hB2BAAB6B5556EAD55532BB6D74C2B9525EB55A47F81555555555555555BABA57),
    .INIT_12(256'h2BE8AB2B55556EA156AAB86D2DACEA874ADC82E9D855AA85555555555506EAA6),
    .INIT_13(256'h3ACBF8BA555555B987EAB86824139DB43EA0E93FBFABAF815AC555555AAABAEB),
    .INIT_14(256'hDEB8AE9E95555550FF7AF9B5C108281CF9F649EA54EFE1455FD6EAAABAAAAAFB),
    .INIT_15(256'hF2EA6ECAD5555541183BA8E5E5AB7918ACE6552011BFDB95404011FABFFEBFFA),
    .INIT_16(256'hF4AA6A5695555414A52BAC82255155592105555555453229555540C5BABFFFFF),
    .INIT_17(256'hFEEEEA46A5555565F57BAD975555555405555555555556319555554551EAAFFF),
    .INIT_18(256'hFCFAAEC5B555567A258BAAD795555555555555555555510AD95555405103AAFB),
    .INIT_19(256'hFF9AFAA5A55556E6169BBE8915555555555555555555562A2C55555555478EAA),
    .INIT_1A(256'hFFABFEA561555D01568BEA5C55555555555555555555546D915555555554293A),
    .INIT_1B(256'hFFF3FFE57955461554EAEA5A55555555555555555555558B61555555555545A6),
    .INIT_1C(256'hFFEBABE94955B89554BAAB3155555555555555555555568CF25555555555550E),
    .INIT_1D(256'h7FF7FFE95555E1D555FA6A615555555555555555555554951885555555555550),
    .INIT_1E(256'hE6FEEFED555661C555AB6911555555555555555555195B6488C5555555555555),
    .INIT_1F(256'hED2DEEAD5555A58554BA2D055555555555555555555646942125555555555555),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_000000_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n122,addra[14:13]}),
    .dia({open_n126,open_n127,open_n128,open_n129,open_n130,open_n131,open_n132,1'b0,open_n133}),
    .rsta(rsta),
    .doa({open_n148,open_n149,open_n150,open_n151,open_n152,open_n153,open_n154,open_n155,inst_doa_i0_001}));
  // address_offset=0;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFCBFE7FBBEFFFFFFFFFEFEFEBFB92EBBFEEFEFFFFFFFFFFFFFFFFFFFFFFAABE),
    .INIT_01(256'hFFDEAFFEB9AAAAAAAAAADAEFABAF79EBBFEEF7FAAAAAAAAFFFFFFFFFFEE001F4),
    .INIT_02(256'hFFEEEBDFBD7AAAAAAAABDEEFBFB9ACBBBBFB9FFAAAABEFFEFA5557AE907BAFCB),
    .INIT_03(256'hFFEEFAFBEE7AAAAAAAAB6EEFAFB4F87BBBEE6EAFAAAFFB956BEAB906EBFFFD2F),
    .INIT_04(256'hFFEFAFBFAEFAAAAAAAAB2EEEFFE7DF2BBBAC7AAFAABE97EBFFA556FFFEBBF2FF),
    .INIT_05(256'hFFEFBEBEEFBAAAAABFAE3EEEBBC2AA6FFBBCAAAAAAB9AFFFA41BEAFABAAF9BFF),
    .INIT_06(256'hFFEF9FBD6EEAAAAABFAF7BFAFB97F7CFFBFEEAAAAABBFFBC0FEEAFAAABBDBFFF),
    .INIT_07(256'hFFEECBAF3EAAAAAABFADFFBBEF5EBA8FFAFFEAAAAAAFF5DBAFEBEAAAABE2FFFF),
    .INIT_08(256'hFFDECFAB3EAABFAABFF8BABAFE39FE8BFBFBAAAAEFFB5BEFEAFEAAAAAAF517BE),
    .INIT_09(256'hFFDEDBABEEAAABEABFFCEBAAFA6EBEE2FFFAAAAABE96FFFEBFEABEAAAAFFEBE9),
    .INIT_0A(256'hFFCFE7BBEEAAAAFABFB9EBAFEDAF7FB6FFEEAAAFF9BAFFABEAAFFEAAABEFAAAA),
    .INIT_0B(256'hFFCBF3BBBAAABEFEBEB6EB9FEC7EAFB6BFEEAEAFDEFBFAFAAAABFEABEAB8AB55),
    .INIT_0C(256'hFFDFE6FAFAAAAFFBEAB7EBDBBC9FDBF1BFBEAFBEFFFEBFFFFFFFEAAAAAB8FFFF),
    .INIT_0D(256'hFFDFF3FBEFEAEEFEFAF6EFAFB4A2DFF4BFBEAFEFFFFEAAAAAAAAFFAAAAAE7FFF),
    .INIT_0E(256'hFFE7F6FBFBFEBBBFAFF6FFFFF3EAAAE9BEEFBEBFFFFFFFFFFFFFEAFFFAAB9BFF),
    .INIT_0F(256'h7FF3F9EEFFBEBEEAFBE7FE7EE6FDF6E8FEFAEFFFFFFFFFFFFFFFFFEAFEAEFEFF),
    .INIT_10(256'hE7E7B8EEFFEBFFFABFBBFE6ED6BAA2ACFFFEBFFEAFFFFFFFFFFFFFFFEBFFBE2F),
    .INIT_11(256'hFDF2FCFEFFFEBFBFFF9FEFFBD65E04EDFBFFFAF907BFFFFFFFFFFFFFFFAFEFDB),
    .INIT_12(256'hBF76FDBEFFFFEBEFFE9BEFBBC0435179EFE2B9117AFFAAAFFFFFFFFFFFFEBFE5),
    .INIT_13(256'hBFA4EF6FFFFFFFABA90FEFFA8648731AEF5A06914054007BFAEFFFFFFAAAAFBC),
    .INIT_14(256'hEBE1FA7BBFFFFFFA418FAEAF3A874E827954FF45FA001ABFE56EBFFFEFFFFFAF),
    .INIT_15(256'hEBBCFB7BBFFFFFED6F8EFEAE3AD3DEF5111BAAFFEE406ABFFFAAAFAFEAABEAAF),
    .INIT_16(256'hFBFEBFAFFFFFFEBF5A9EFAE9FAAAAAAF9EFAAAAAAABA84ABFFFFFE6BAFEAAAAA),
    .INIT_17(256'hFDBBBFEEEFFFFFEE1ADEFBFDAAAAAAABFAAAAAAAAAAAAC4BBFFFFFFAAFBFFAAA),
    .INIT_18(256'hFF7FFBAFEFFFFED0BA6EFFB9EAAAAAAAAAAAAAAAAAAAAEE57BFFFFEAFEAEFFAE),
    .INIT_19(256'hFF7FAFEFBFFFFD1BEB6EEBA7EAAAAAAAAAAAAAAAAAAAA80507FFFFFFFFF93BFF),
    .INIT_1A(256'hFF8EABFFFBFFF06EAB7EAFF3AAAAAAAAAAAAAAAAAAAAABC7BEFFFFFFFFFEC7EF),
    .INIT_1B(256'hFFDBAABFEBFFE9AAAB2FAFE7AAAAAAAAAAAAAAAAAAAAAAF4ABFFFFFFFFFFEE5A),
    .INIT_1C(256'hFFF2FEBBEBFF97EAAB2FAE9AAAAAAAAAAAAAAAAAAAAAAB6B4EFFFFFFFFFFFFB5),
    .INIT_1D(256'hFFF9EABBFFFF1F2AAA2FEEDEAAAAAAAAAAAAAAAAAAAAAB2AE2AFFFFFFFFFFFFB),
    .INIT_1E(256'h5BFCBABBFFFC503AAA7EEFFEAAAAAAAAAAAAAAAAAAEEACFB142FFFFFFFFFFFFF),
    .INIT_1F(256'hE5BE7BFBFFFF96FAAA7EEBAAAAAAAAAAAAAAAAAAAA9BBCFFC20FFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_000000_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n181,addra[14:13]}),
    .dia({open_n185,open_n186,open_n187,open_n188,open_n189,open_n190,open_n191,1'b0,open_n192}),
    .rsta(rsta),
    .doa({open_n207,open_n208,open_n209,open_n210,open_n211,open_n212,open_n213,open_n214,inst_doa_i0_002}));
  // address_offset=0;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFD7FFDCB09FFFFFFFFF41F00FFF877FC3FF289FFFFFFFFFFFFFFFFFFF7D5FDD),
    .INIT_01(256'hFFDD5D2F973555555557F7D827D42B5F61D78E7D5555555F575555555D25D535),
    .INIT_02(256'hFF45D7FD35F755555557B5DAA57CB3FFEDF4D1775557DDDF2A75550A95D0D791),
    .INIT_03(256'hFF45F5CB94F55555555567F29557AE5F6FF3455F555F5C3D401F4B7CBF57DD7F),
    .INIT_04(256'hFF675F773F9555555555FDD095F0B0DDE7DAD55F557F9DB5FDC5DCBDFF77CEFF),
    .INIT_05(256'hFF67C57ABD7555557F5DFFF8F57561652762F55555773F5DED5A95F5755D1FFF),
    .INIT_06(256'hFF477F775DD555557F565FE0F76C06BF2D29DD55557757C754195F55577FBFFF),
    .INIT_07(256'hFF65DF540D5555557F559F60FD72CA712D89D555557DCF787097FD5557D67FFF),
    .INIT_08(256'hFFFD515565557F557FF7F7EBF5CD02F10C0F5555DF7C7AB2BFFFFD5555CD7D21),
    .INIT_09(256'hFFFD5955A5555FD57FF35F61F6F0200F02255555553CA2A15DFD555555F5D429),
    .INIT_0A(256'hFF7F4777DD5557F77F5B7F41D930C2A90ABD555DC32D28D7FFF5555557DD7DFD),
    .INIT_0B(256'hFF5FE5F7FF555FBDFF5457D35B4308AAE81D5FF513042DFD75555555557FA1D5),
    .INIT_0C(256'hFFF3F3F7F5557F8F5F54D7B7C3301C8DE87D5FF52201FFFFFFFFD5555577BFFF),
    .INIT_0D(256'hFFD1F4549FD5FBEBF5D5D7AFE64B10A760FD55580021D55557DDFFF7555DEFFF),
    .INIT_0E(256'hFFCDD65685FF7EF2FFF5DF658630E30A415F7FC8A802828002A89F7FF55753FF),
    .INIT_0F(256'h6FCDD3D7AAFD7DB52555FD6D0F012F0181F5D08AA02A0000000AA8357F55F6FF),
    .INIT_10(256'hEDF3F7DF0017D58542497D5D958C344B03D74A2B5802020A800000AA1DFF74DF),
    .INIT_11(256'h7975FF3D0003FFCA80F35C5438C37E0987D8270974400000000000A0A2FFFD2B),
    .INIT_12(256'h14F4773F020A15DAA3F7FC9416F47F4B376DEB74670A7DD0AAA002AA8AA97F59),
    .INIT_13(256'h85C5747D82AA827ED957D6B7B029D7D0175676A57D7F5D448F300000AD7F5F7F),
    .INIT_14(256'hEFD6FFC7E02A808FFDBDD45060A4308E7E31E9BDF87DF8A00DC1D55557FFFFDD),
    .INIT_15(256'hDB7F9FEFE002801AA8955E58CABE621EDE502A000077ED682220A8DFFFFDD57F),
    .INIT_16(256'hF25715A9400001E2701756F5CAA2A221388AAAAAAA0A993E00008AC2DFDD5555),
    .INIT_17(256'hF7F77723D8002AB8E05754C2AAA828A2AAAAAAAAAAAAA53A480000A8027F5555),
    .INIT_18(256'hFEDFD74058002335284777482AAAAAA2AAAAAAAAAAAAA8256C0008150029DD5D),
    .INIT_19(256'hFF675FDAD80003D2A845757D2AAAAAAAAAAAAAAAAA82A19D540000000009A5FF),
    .INIT_1A(256'hFF7F5FD03E0026AAAACF5D8CAAAAAAAAAAAAAAAAAAAAA256CA80000020032F1F),
    .INIT_1B(256'hFFD97DDAB6001B2AAADFFF24AAAAAAAAAAAAAAAAAAAAA00D34000000280030F9),
    .INIT_1C(256'hFFD7FD7E9600D6AAAAFFFF58AAAAAAAAAAAAAAAAAAAAAAE0D9000000000000CD),
    .INIT_1D(256'h3FF3D576A8025BEAA8DFBD9AAAAAAAAAAAAAAAAAAAAAAAC0845000000000000E),
    .INIT_1E(256'h5BF7F576A009184AAA7D9E32AAAAAAAAAAAAAAAAAAC2A3C2E4F0000000000000),
    .INIT_1F(256'h763E77FEA00A700AAA5F9E02AAAAAAAAAAAAAAAAAA80251CB6D8000000000008),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_000000_003 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n240,addra[14:13]}),
    .dia({open_n244,open_n245,open_n246,open_n247,open_n248,open_n249,open_n250,1'b0,open_n251}),
    .rsta(rsta),
    .doa({open_n266,open_n267,open_n268,open_n269,open_n270,open_n271,open_n272,open_n273,inst_doa_i0_003}));
  // address_offset=0;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFF65573FF57555555555F77F5557E1D5FD57DD75555555555555555555FF75FF),
    .INIT_01(256'hFF65575FFEF55555555565777D5FB4D5DD5771D555555555FFFFFFFFF7D22052),
    .INIT_02(256'hFF5D55675E9555555555ED75F55EFC555D5FC755555557F75D2AA8D76005DFC7),
    .INIT_03(256'hFF7D557F5F35555555573D5F75725FB55D7F3D555555FFE2377FF4AB5DFD769F),
    .INIT_04(256'hFF7D5551757555555557955D555B4F35D55F35555557E057FF522BDF5555DBFF),
    .INIT_05(256'hFF7DDD5F755555555557957555E9D59DD5DFD555555E57FF70075D555557CFFF),
    .INIT_06(256'hFF7D655EB5555555555D357F5561F967D5D755555555FDF281FDD55555567FFF),
    .INIT_07(256'hFF5D4D5D95555555555E75775587FD45D57D555555577825FFF555555571FFFF),
    .INIT_08(256'hFF65C7579D5555555554D5DD551E7FE5FFF5555555D585FD77555555555208D7),
    .INIT_09(256'hFF45EF57FD5555555556D5F55FBF7F53FDF555557F6B7D5DD5555555555F5DF4),
    .INIT_0A(256'hFFE5FB5575555755557ED5D55E7F3D51F555555556DFD7F55555555555577FFF),
    .INIT_0B(256'hFFED7B55555555D55571D5655C3F7F51D7D5555767FFF5555555555555547CAA),
    .INIT_0C(256'hFFC57355555575FD557955E5F6CF6FD0D7555557FDFDD555555555555556FFFF),
    .INIT_0D(256'hFFC759D7D5557F75557B55D57B7FE7785FD5557FFFDD5555557D555555553FFF),
    .INIT_0E(256'h7FDB7BD77555557DF559551DF9F7D7F67D5557F757FD7D7FFD57D755555567FF),
    .INIT_0F(256'hBFDB74D757D55577D5FB5597FBFED3FCFF5557755FD5FFFFFFF557F7555551FF),
    .INIT_10(256'h5BF15E55FFD555FFFF7F5795C3DD797CF55DF5FF75FDFDF57FFFFF55DD555FBF),
    .INIT_11(256'hF6715657FFFDD5F57FED5537C18522FE7D7FDFD683FFFFFFFFFFFF5F5F7557EF),
    .INIT_12(256'hFD9BDE57FDF5DD755FED57FF4A81A01475D3D40297FF7DFF555FFD55755F55F8),
    .INIT_13(256'h5FF8DFB5FD557F7DFE855DD741060AAD7D0FABC0A882023F7FFFFFFFFD55D556),
    .INIT_14(256'hFD5857155FD57F7F2A455DDF1F4185CBB62034828FA08D7FF2BDD55555555557),
    .INIT_15(256'hF554F595DFFD7FF615ED57771F41274822057F5557A8BD57D7D575D555555555),
    .INIT_16(256'hFDDD77FD7FFFFF5F2DED577C9FF7DFF4EFDFFFFFFF5D607DFFFF5D9755555555),
    .INIT_17(256'hFCD5555D57FFD57FAD0D557C7FFFFFFFFFFFFFFFFFFFD0A777FFFF7FF7D55555),
    .INIT_18(256'hFDB5555F77FFDFE87DBD55F67FFFFFFFFFFFFFFFFFFFFD789FFFF7FFF7577555),
    .INIT_19(256'hFF3D555557FFF487FD1D75707FFFFFFFFFFFFFFFFFFFFCA089FFFFFFFFD6DF55),
    .INIT_1A(256'hFFC5555FFDFFDA97FFB575FBFFFFFFFFFFFFFFFFFFFFFF09FD7FFFFFDFFF72D5),
    .INIT_1B(256'hFFE7555D55FFDEFFFFB5D7F1FFFFFFFFFFFFFFFFFFFFFF707FFFFFFFD7FFFF0F),
    .INIT_1C(256'hFFD3555D75FFC37FFF3555CDFFFFFFFFFFFFFFFFFFFFFFB705FFFFFFFFFFFFD8),
    .INIT_1D(256'h7FFED5555FFDA43FFF15D54FFFFFFFFFFFFFFFFFFFFFFD3FD97FFFFFFFFFFFFD),
    .INIT_1E(256'h0DFCD55D5FF4883FFD955767FFFFFFFFFFFFFFFFFF97F61F203FFFFFFFFFFFFF),
    .INIT_1F(256'hDA5F355D5FF5417FFFB75FF7FFFFFFFFFFFFFFFFFFE5F0616387FFFFFFFFFFF7),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_000000_004 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n299,addra[14:13]}),
    .dia({open_n303,open_n304,open_n305,open_n306,open_n307,open_n308,open_n309,1'b0,open_n310}),
    .rsta(rsta),
    .doa({open_n325,open_n326,open_n327,open_n328,open_n329,open_n330,open_n331,open_n332,inst_doa_i0_004}));
  // address_offset=0;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFDAF9BF7ADBBFFFFFFF8E8E83AA31FE3BA8ACBFFFFFFFFFEFFABAFFFEBF8138),
    .INIT_01(256'hFFFAFEED631FBFFFFFFBBBCA02EBE3EA6ABEEEBAFFFFFEAEFBAFFEBAACDD1934),
    .INIT_02(256'hFFDEEFEBAFEFBFFFFFFABA8ABFE2682E6FE2FEFAFFEFFBFC757FA8696A897B97),
    .INIT_03(256'hFFDAFBF3F8FFFFFFFFFA5B9D0BEDEBFE7FDFCFAAFFFEA62B1F01634C83FEFE5F),
    .INIT_04(256'hFFDBFFB289EFFFFFFFFF4A8CFFCBFB1BA7CABFFAFFF87CDEFF27A8FBBEBBC1BB),
    .INIT_05(256'hFFDB3EFD9FBFFFFFFFF97FAC7F95C5CFA22F6BFFFFE2DAEE0D7482BFBEAE63FF),
    .INIT_06(256'hFFCBFBFBCBFFFFFFFFFE7FF1BA3AAF8CA7BDFFFFFFFBAB6162FD7BFFFFBA6FFF),
    .INIT_07(256'hFFCAA2FC5FFFFFFFFFFABFF6FFFAE543B0FABFFFFFEBAA26FA8BFFFFFF94AFFF),
    .INIT_08(256'hFFAAA7FE3AFFFFBFFFF87B39BC3EBA97ABA6FFFFFEA7B3FBB5BEFFFFFFDBF861),
    .INIT_09(256'hFFEBF6FB8AFFEEFFFFE0AF53A1293890FFFFFFFFF8BCBBAD3BEABFFFFFFFB0C5),
    .INIT_0A(256'hFFCF8FBB8FFFF8BFFFF3BE1EAF2EFE29FF8AFFFE876EEB9AEFEBFFFFFFFA8554),
    .INIT_0B(256'hFFC6B7BFEBFFF8AAEAA7AF23D8EF4E2DFFEAFAFBFBBEA3EFFEFBEFFFFFE510BA),
    .INIT_0C(256'hFFF3C0F9AAFFCAF6EAEDBEFE787EAE22BE6FFFEDAFFD2EAAAAABEBFFFFF9BFFF),
    .INIT_0D(256'hEBFEE4FBABFFDDA9ABF8AE0E6F5FBADD7B3FEBDFFFF941554402EBFBFFFABFFF),
    .INIT_0E(256'hBBCBE9BAB2BFA34BCAFAEF2BA3B593D73CFFF8EFFFEAAAAAAAAAD1FAFFFEABFB),
    .INIT_0F(256'hEFF6FAFAFB7EFCF7E7DAFF9DC6ABEB90F9BFA7BFFFFFEFFFFFFFAAF1EBFEA0FF),
    .INIT_10(256'h8ED7E1A8BE9FFEEFAAE6FDA8F92F6454F3EB7FEE3BFFFFFFFFFEEBAAD3FFF80E),
    .INIT_11(256'hEAB0F869FAE86A6EFFEBE92EACE80C80F3FABAA359FFFFFFFFFFFFFFEB1AFEB3),
    .INIT_12(256'h6CEDFA29FABEC7DAAEC2AA32C55EF6B3FE93E3F6B7FB3DAFFFFFFFFFFAE9FF8A),
    .INIT_13(256'h4F1BFFDBBBFFEA5FA20FBFA743A8A8708AEF464886FC51CBFABBEBAFF9412FE8),
    .INIT_14(256'h96B3BDDB2FFFFFAFC9AFFF7A9894F9F6F337CE203BCB381F8FC96EFFFEFABFEE),
    .INIT_15(256'hC7ACBFA72FFFFFBEEFBBFCD9B18B99FA7FD2D5EFE97F887FF9401D7AAFBFEFFF),
    .INIT_16(256'hF3ACEA0FBFFFFBF9F6FAF8BF2551154A9171555555F0ED3ABAAAB59A7AFFFFFF),
    .INIT_17(256'hFA6FFA49DBFFFFED429AF9F8554145555555555555551E926FFFFAC11B6EFFFF),
    .INIT_18(256'hFFBFEB9B9BFFFAF3C75AFF7595555555555555555555545EFAFFFFFEE85DEBBF),
    .INIT_19(256'hFFABFFCA3BFFEE10563ADB7ED5555555555555555555575B8ABFFFFFEAA7E2BF),
    .INIT_1A(256'hFB5FFFEF8BFFF5BC54EFDBA55555555555555555555550BBB5EFFFFFFFFABEFA),
    .INIT_1B(256'hFFE6FFFB86FFD684558B49925555555555555555555554C66EEFFFFFFFFFF9F1),
    .INIT_1C(256'hEFF4BFFBF2FE95C554CF089F55555555555555555555543D68BFFFFFFFFFFEBA),
    .INIT_1D(256'h7FF6EFF2FFFB275555AFCDC05555555555555555555550D0407FFFFFFFFFFFFF),
    .INIT_1E(256'h67F96FF2FFEDE70555EE8F8D555555555555555554085AE4B87BFFFFFFFFFFFF),
    .INIT_1F(256'hDA2D7BF7FFFE649557E98679555555555555555551921EFF14CEFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_000000_005 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n358,addra[14:13]}),
    .dia({open_n362,open_n363,open_n364,open_n365,open_n366,open_n367,open_n368,1'b0,open_n369}),
    .rsta(rsta),
    .doa({open_n384,open_n385,open_n386,open_n387,open_n388,open_n389,open_n390,open_n391,inst_doa_i0_005}));
  // address_offset=0;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFEBAFED703EEAAAAAAA82E14FFF4BEB86FE547AAAAAAAAABAAFEFAAABABAEFE),
    .INIT_01(256'hFFAEAA1F2A2AAAAAAAAAFAB15FA817AB86A81DAAAAAAAAABFAAFFEBAAA4BF9B6),
    .INIT_02(256'hFF8EAABE3EBAAAAAAAAB7AE09ABC47FBC6B862AAAAAAAFBAC06FF8442AC3AB62),
    .INIT_03(256'hFF9AAAC768AAAAAAAAAA5AF12EBB43AB96B18AAAAAABA86F55AEC6E86EFFBABF),
    .INIT_04(256'hFF8ABAB33E2AAAAAAAABBEF16AF064EE0AA7EAAAAAAF782FBFC7ED2BEAAAACFF),
    .INIT_05(256'hFF8ACEB46AAAAAAAAAAFBAC4EABA429A4F83FAAAAABB7EEBDAA42AEAAAAA2FFF),
    .INIT_06(256'hFF8AEEAAEEAAAAAAAAAD6A94AB99597E4E46EAAAAAAAAA83E016AEAAAABF7FFF),
    .INIT_07(256'hFF9AEFAE7EAAAAAAAAAA7AD0AAB655BA1B06EAAAAAAFCF35552AAAAAAAF9BFFF),
    .INIT_08(256'hFFFEAFAA8AAAAAAAAAABAADBEA874632004FAAAAABBCA5541FEAAAAAAAFEBC1A),
    .INIT_09(256'hFFFEA2AB5AAAABAAAABBAA96F984150F400EAAAABA3C1402EEAAAAAAAABBFA51),
    .INIT_0A(256'hFFFA8EAAEAAAABEAAAB6AB83E640C017003EAAAAE305002BAAAAAAAAAAAEBAAA),
    .INIT_0B(256'hFFABCFAABAAAAF3EAAA4AAEAA7911505402EAAAB25401FBAAAAAAAAAAABF40EA),
    .INIT_0C(256'hFFEBBBABFAAABF4FAAAAEB2FC331751B00BAAABA1002FFFFFFFEAAAAAAAB7FFF),
    .INIT_0D(256'hFFE2BFE86EAAA7D3FABAEB5FDB8D655B84EAAAA40007FEAAABEEBEAAAAAEDFFF),
    .INIT_0E(256'hFFCEA8A90EEABDE57FAAAA1A5D50150582AAAF400014000000006BAFAAABA3FF),
    .INIT_0F(256'hDFCAB3AC00AAAA580AFAABAE1C56194642EAE800000000000000001EBEAAF1FF),
    .INIT_10(256'hCAEEBAEF002EAA0001C2ABAF6F4119870AAEC01491000000000114002EAAA8EF),
    .INIT_11(256'hE3BAEFFE0503FFC10073AE2964D7BC570AA40002FD0000000000000001FFAA07),
    .INIT_12(256'h6EBDAB3F05402AE1542BAC6838ADBB825B9912F899058210000000000047EAA6),
    .INIT_13(256'h6FDFACEE440001B016AAAC693C07DDE56BA6E56DFBABAE941014005552BEAABF),
    .INIT_14(256'hDFF8EABBC0000005ED6EACE5F6422A4EBCAF79E111ABF9004ED2EAAAABAFEAAA),
    .INIT_15(256'hE7BB7B9FC00000014B2AA8E4EE8F7AD8B98EEAEFFF6AD380111057AFFAAAAAAA),
    .INIT_16(256'hF5AF6A56D0000005BB3AA8D62AAAFAB95EFEAAAAAAFE2241455505C1FFAAAAAA),
    .INIT_17(256'hFBFAEBD7E0000004BB5AAB82EABEBAABFAAAAAAAAAAAF2659000054400BFAAAA),
    .INIT_18(256'hFDEAAAC4E000043E2B5AAB86AAAAAAAAAAAAAAAAAAAAAEDE910000010016EEAA),
    .INIT_19(256'hFF9AAAA0A00016CEEA1AAA99EAAAAAAAAAAAAAAAAAAAAB6E6D4000000556DEEA),
    .INIT_1A(256'hFFFEAAA06400191EAACEFE4AAAAAAAAAAAAAAAAAAAAAAF690510000000053E3F),
    .INIT_1B(256'hFFE6AAA42800337AABEEBF42AAAAAAAAAAAAAAAAAAAAABB705000000000014E6),
    .INIT_1C(256'hFFEBEAA01C0113AAABFAFE57AAAAAAAAAAAAAAAAAAAAAA5B360000000000014F),
    .INIT_1D(256'hFFF3AAAC0405B96AAAAA7E1EAAAAAAAAAAAAAAAAAAFAAFEFFC80000000000005),
    .INIT_1E(256'h67FBBAA80012247AABBA391EAAAAAAAAAAAAAAAAAB3AAA6FC9D4000000000000),
    .INIT_1F(256'hB93D6AAC0000BAAAA9AE3D5EAAAAAAAAAAAAAAAAAA3EB2C3ED61000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_000000_006 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n417,addra[14:13]}),
    .dia({open_n421,open_n422,open_n423,open_n424,open_n425,open_n426,open_n427,1'b0,open_n428}),
    .rsta(rsta),
    .doa({open_n443,open_n444,open_n445,open_n446,open_n447,open_n448,open_n449,open_n450,inst_doa_i0_006}));
  // address_offset=0;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFF9AAB3EFAAAAAAAAAAAFBAFAAABD2AABEAAFEAAAAAAAAAAAAAAAAAAAAFEBAEF),
    .INIT_01(256'hFF9AABAFFDFAAAAAAAAA9ABFBEAF78EAFEAAF2EAAAAAAAAAAFFAABEFFBA003AD),
    .INIT_02(256'hFFAAAA9BA96AAAAAAAAADEBF3AADECAABEAFCBAAAAAAAAEBEED006AB902BEFCB),
    .INIT_03(256'hFFAEAABFAF3AAAAAAAABFEAFFAB1B97AAEBF3EAAAAAAFF90EEBFB817AEAAA96F),
    .INIT_04(256'hFFBEBAAABABAAAAAAAAA6AAEAAA79F3ABAAD3AAAAAABC2AEFEAC16EEAAAAE7FF),
    .INIT_05(256'hFFBEEAAFBAAAAAAAAAAA6AAAAAD6FA6EFAFDEAAAAAADEBBEB00AEEAAAAABCFFF),
    .INIT_06(256'hFFBEDAAD3AAAAAAAAAAAFABFAA96F69AFAFBAAAAAAAAFEF90AFEEAAAAAA9BFFF),
    .INIT_07(256'hFFAE8EAA3AAAAAAAAAADAAFBAA48FE8AEEFEAAAAAAAAB49AFFBAAAAAAAA2FFFF),
    .INIT_08(256'hFF9ACEAB6EAAAAAAAAA8EAE2AA6DBC9AFBFAAAAAAAEA4AFFFBAAAAAAAAB106EB),
    .INIT_09(256'hFF8ADFAAFEAAAAAAAAA9EAFAAF2FBFA3BFFEAAAAAF97FFFEEAAAAAAAAAAEBEBB),
    .INIT_0A(256'hFF9AF3AABAAAABAAAAADEAEAADAF3FE3FFEAAAAAA9FFFFBAAAAAAAAAAAABBFFF),
    .INIT_0B(256'hFFDEB2AAAAAAAAAAAABEEA9AAC3FBFF2FFEAAAAA9BFFFBAAAAAAAAAAAAA8BE55),
    .INIT_0C(256'hFFCAB3AAAAAABAFEAAB6AADEF9CF9FA4BFAAAAABFFFEEAAAAAAAAAAAAAA9FFFF),
    .INIT_0D(256'hFFCBA3ABEAAABFBEAAA7AAEAB5B7DBB4BFEAAABFFFFEAAAAAABEAAAAAAAA3FFF),
    .INIT_0E(256'hBFE7B7EBFAAAAAAEFAA6AAAEF6FBABF9BEAAABFFFFFFFFFFFFFFEFAAAAAA9BFF),
    .INIT_0F(256'h3FE7A8EAFFEAAABBFAA7AB6BF6FDE7FCFFAAABFFFFFFFFFFFFFFFFFBAAAAAAFF),
    .INIT_10(256'hA7F6ADAAFFEEAAFFFFFFAA6AC2FBA6BCFAAABFFEBEFFFFFFFFFFFFFFEEAAAF7F),
    .INIT_11(256'hB8B2A9EBFFFEEAFFFFDEAABBD24A10FDFEBFFAED03FFFFFFFFFFFFFFFFBAABDF),
    .INIT_12(256'hBA62EDABFFFFEEBFFE8EABFF8506402DBAE7A8416BFFAABFFFFFFFFFFFBEEAF4),
    .INIT_13(256'hAAE1EB3AFFFFFFBBBD4AAAFB870D261EBE0C1E871501013FFABFFFFFFAAAEAA9),
    .INIT_14(256'hFEB4AB3ABFFFFFFF13CAABAF7FCF1AD47914BA1FAB1142EFF17EEAAAAAAAAAAB),
    .INIT_15(256'hFAA8EA6AFFFFFFF92B8EABFF6FB68BE4007AFFEFFEC07ABFEBEABBEAAAAAAAAA),
    .INIT_16(256'hFEEAFBFEBFFFFFFF0FCEABBCAFFBEFFAFFFFFFFFFFFFC0ABFFFFEE6BBAAAAAAA),
    .INIT_17(256'hFCEAEAEEAFFFFFEF4FBEABBCBFFFFFFFFFFFFFFFFFFFE91BBFFFFFAFFBEAAAAA),
    .INIT_18(256'hFE7AAAEFBFFFFED1EFEEAAF8BFFFFFFFFFFFFFFFFFFFFFA06BFFFFFFFBABBAAA),
    .INIT_19(256'hFF3EAAAFEFFFF97AFEFEBAB2FFFFFFFFFFFFFFFFFFFFFC0046FFFFFFFFE96FAA),
    .INIT_1A(256'hFF8AAAAFEFFFE56FFE3AEAF7FFFFFFFFFFFFFFFFFFFFFF96BEFFFFFFFFFF90FA),
    .INIT_1B(256'hFFDBAAAFFBFFFCFFFF3AEBFEFFFFFFFFFFFFFFFFFFFFFFBDAFFFFFFFFFFFFF0F),
    .INIT_1C(256'hFFE3AAABFBFFBFBFFF7AABFFFFFFFFFFFFFFFFFFFFFFFEFBDAFFFFFFFFFFFFE4),
    .INIT_1D(256'hFFFDEAABFFFE4EBFFF2AEAFFFFFFFFFFFFFFFFFFFFFFFE3FE2BFFFFFFFFFFFFE),
    .INIT_1E(256'hCEFCEAAFFFFC41BFFE2AEBAFFFFFFFFFFFFFFFFFFFABF8AB503FFFFFFFFFFFFF),
    .INIT_1F(256'hE5AFFAAFFFFF87BFFF3BEFBFFFFFFFFFFFFFFFFFFF9AF9BBD74FFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_000000_007 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n476,addra[14:13]}),
    .dia({open_n480,open_n481,open_n482,open_n483,open_n484,open_n485,open_n486,1'b0,open_n487}),
    .rsta(rsta),
    .doa({open_n502,open_n503,open_n504,open_n505,open_n506,open_n507,open_n508,open_n509,inst_doa_i0_007}));
  // address_offset=8192;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hEDBFB9ABFFFEAFAFFDA8D6BBFFFFFFFFFFFFFFFFEADA2A9BCD13FFFFFFFFFFFF),
    .INIT_01(256'hBEDAB869BFFCC6BEB9F887AFFFFFFFFFFFFFFFFFEE2B049BA61BFFFFFFFFFFFF),
    .INIT_02(256'hFFAC2928BFFF9EBEBB7BB96FFFFFFFFFFFFFFFFFEF73D19EBD4FFFFFFFFFFFCF),
    .INIT_03(256'hFFAECADCBFFADEBEB3E6FA3FFFFFFFFFFFFFFFFFEBF37EAEBB9AFAFFFFFFFE25),
    .INIT_04(256'h0AAAEE6DBFC59FFEB0E248EFFFFFFFFFFFFFFFFFEAF3747AEA147AFFFFFFFFD5),
    .INIT_05(256'hE6A6BE66FFFE3FEEB9B7CFAFFFFFFFFFFFFFFFFFEAF1FAEBEAA99FFFFFFFFF8A),
    .INIT_06(256'hDBAEAFBA2F68BFFFA863F42FFFFFFFFFFFFFFFFFEAF356FEEAE4F3FFFFFFFFB8),
    .INIT_07(256'hF8E6BF9C6EA6EBFBEC6F6C7FFFFFFFFFFFFFFFFFFFEDC6FBABA0F6FFFFBC3FFF),
    .INIT_08(256'hFFBD1B8A3FE6BEAFECAE748BFFFFFFFFFFFFFFFFFFEFEBBBA3F9BBFFFFF6E3FF),
    .INIT_09(256'hFE9B06EEBE26BFFFFCDBF90EFFFFFFFFFFFFFFFFFFEF5FB8304EBEFFFFFE6A7F),
    .INIT_0A(256'hFF9E4CA6FE7FFFEAF28CCA1FFFFFFFFFFFFFFFFFFFEFAF5DAFE2CDFFFFFE39F6),
    .INIT_0B(256'hFEEB9C32BE0BFCE4A6DF4524AFFFFFFFFFFFFFFFFFEFF933BABE727FFFFAC3D4),
    .INIT_0C(256'hFFFEFB5FF20FBBB4F4D95EDAABFFFFFFFFFFFFFFFFFFE69AEFFFED6FFFFFF1FB),
    .INIT_0D(256'hFFF4BBE5FB4FB0AAE9D8370F6ABFFFFFFFFFFFFFFFFADEEFFFFFE0EFFFFFE97E),
    .INIT_0E(256'hFFF96E3DFB7EDC1A0700F2AB5BBFFFFFFFFFFFFFFFFA838AFFEBC5FFFFFFEE1F),
    .INIT_0F(256'hFFFFA2EFFDAF4001804DCF6EEFBFFFFFFFFFFFFFFEEF1B6AFFEBB89FFFFFFEFF),
    .INIT_10(256'hFFFFDE757DAF5169C1CAC4E2B3BFFFFFFFFFFFFFFEB833AABFEBA47BBFFFFF97),
    .INIT_11(256'hFFFF4E8D99AB003EF6DDB344E0FFEFFFFFFFFFFFEA35FBBFFFEBEFABFFFFFFC4),
    .INIT_12(256'hFFFFD1E248BA02EA82BB0864DAEFFBBFFFFFFFFFE816BBFFFFFFEBCBFFFFFFF6),
    .INIT_13(256'hFFFFECD4E73B13AFF2D41255666AFBBFFFFFFFFEA51EFFEABFFFEF16FFFFFFFC),
    .INIT_14(256'hFFFFF47B0E6B5FFFF34BAC245E2AFFABFAFFFFFE9B6EEFFAFAFBFD2FFFFFFFFF),
    .INIT_15(256'hFFFFFDBC006F67FFF62DA0819E7EBEFFFFFFFFFB6CC3EAAAFEEBFF3BFFFFFFFF),
    .INIT_16(256'hFFFFFE23BDAF6BFFFB26FF38FA72BAABFEFFFFEE96DFF0B1BBABFFB3FFFFFFFF),
    .INIT_17(256'hFFFFFF6F54BA2FFFF8CDFFF255EAB5AEBABFEFBA4CA5EFFEA05FAFDAAEAFFFFF),
    .INIT_18(256'hFFFFFFF90A3B03FFFD5BFF9F28C5B8EEEFBFEAB5E53D142907EBAF18DFFFFFFF),
    .INIT_19(256'hFFFFFFD4EF4F17FFFFAFFCC3EA373EEE9ABFFACC8DD00007397EBF2583AFFFFF),
    .INIT_1A(256'hFFFFFFF461DF07FFFC4FFC3DFE4DF6AFB3AFF9368000691D03DBBFA0C71FFFFF),
    .INIT_1B(256'hFFFFFFD1AADE13FFFEAFFFFEFC0939AFCFEEB2300C8EFFFF2C32EABD47FFFFFF),
    .INIT_1C(256'hFFFFFFC3123AAFFFFEFFF7FBBF4AD0FFDFAB078C3013AAAAED41EAB2892FFFFF),
    .INIT_1D(256'hFFFFFFD10CFAAFFFFF5FF52DFF3BD2FF66AFE7111FFFFAAD7B4AEF62AF8BFFFF),
    .INIT_1E(256'hFFFFFFD25A2E93FFFFAFF165BFA966AB62EFB52B67FFFFFFEA17FFFBDFCBFFFF),
    .INIT_1F(256'hFFFFFFEE47FEEFFFFF6FF211BFD7F2AAE34A38F3A7FFFFFFF51BFA8A4B0BFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_008192_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n535,addra[14:13]}),
    .dia({open_n539,open_n540,open_n541,open_n542,open_n543,open_n544,open_n545,1'b0,open_n546}),
    .rsta(rsta),
    .doa({open_n561,open_n562,open_n563,open_n564,open_n565,open_n566,open_n567,open_n568,inst_doa_i1_000}));
  // address_offset=8192;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hEA8FBBA95554C15555BA29D5555555555555555554D1D0212FC5555555555555),
    .INIT_01(256'hBEA94FEB5556995551EA68855555555555555555543427915AE1555555555555),
    .INIT_02(256'hBFAAEFAA5554A55552295005555555555555555555B0DCE55675555555555565),
    .INIT_03(256'h2FAEBA7B555265555B7D52155555555555555555554997455528555555555420),
    .INIT_04(256'h2AAAEE9B556155555B3D435555555555555555555543919555A3955555555564),
    .INIT_05(256'hBEAABEDA555A95555269D3155555555555555555555A5C555502E5555555552E),
    .INIT_06(256'hEEA5AF9695B3155552A981955555555555555555555A40555546F95555555511),
    .INIT_07(256'hF0AA6FA2946C555556E5CA955555555555555555555480550159F45555569555),
    .INIT_08(256'hFE6BFBB59570555556A5D8A555555555555555555554D1415456B5555555D955),
    .INIT_09(256'hFEBA7AE55469555553B4820555555555555555555554A557311090555555ED95),
    .INIT_0A(256'hFF5A8BA954C5554052F5CAD555555555555555555554C58C8545165555558388),
    .INIT_0B(256'hFFF688ED146554B043E726F65555555555555555555556261555B39555502F3C),
    .INIT_0C(256'hFFFE8B795BA55545E9E3657D155555555555555555555B8C5555464555554AF1),
    .INIT_0D(256'hFFF1FFCE51A55A005C66789A955555555555555555556BE155554B05555542BF),
    .INIT_0E(256'hFFFFE67652554D04B736ED4B6455555555555555555533A555556855555554FF),
    .INIT_0F(256'hFFFCF8955755A0003C7BAC83845555555555555555559E95555554E55555542B),
    .INIT_10(256'hFFFFFD7A9215A23A002AB68FED555555555555555556215555555A515555551E),
    .INIT_11(256'hFFFFB90BE215A1944F268D27B255555555555555558CD0555555541155555563),
    .INIT_12(256'hFFFFC649E705A05567561E9B885555555555555556271555555555015555555A),
    .INIT_13(256'hFFFFFA474385B6FFFB5FD069C79555555555555559D841555555557955555556),
    .INIT_14(256'hFFFFF8AC9695B3FFFD8D4413AB055455555555556F751555555556C555555555),
    .INIT_15(256'hFFFFFD2BAA959BFFFDFFE8023CC5575555555555A9F940005555553555555555),
    .INIT_16(256'hFFFFFF2013159BFFF9A3FEB0576D53155555555481B00EF10505556955555555),
    .INIT_17(256'hFFFFFF907B559FFFFF31FFFF442454155555555343F115500115556144055555),
    .INIT_18(256'hFFFFFFE2A215B3FFFD3AFFAFB2AA58555D555519EFC41412F92555A4A5155555),
    .INIT_19(256'hFFFFFFD41225B3FFFDEFFFD7E552995508555420DF400001A69555B5AC455555),
    .INIT_1A(256'hFFFFFFF4ADA5A3FFFFCFFC32FB2A5855215550DD0002EBE000A15521B6E55555),
    .INIT_1B(256'hFFFFFFD5D1E5A3FFFE4FFB3CFF43DE556555539006D155546000552C49555555),
    .INIT_1C(256'hFFFFFFC769C53FFFFF1FFF3DFF93A6552155D1030BE95555454A5527A6855555),
    .INIT_1D(256'hFFFFFFC111852FFFFFBFF97DBF0690557954C5DBBFFFFFFB840455E356D15555),
    .INIT_1E(256'hFFFFFFC349C51BFFFFAFF91DFF8DA455294629AA3BFFFFFFE63955626E915555),
    .INIT_1F(256'hFFFFFFF3435552FFFFBFFB41FFEEE054A98DA3F2E3FFFFFFFE11551280515555),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_008192_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n594,addra[14:13]}),
    .dia({open_n598,open_n599,open_n600,open_n601,open_n602,open_n603,open_n604,1'b0,open_n605}),
    .rsta(rsta),
    .doa({open_n620,open_n621,open_n622,open_n623,open_n624,open_n625,open_n626,open_n627,inst_doa_i1_001}));
  // address_offset=8192;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hBE566EFFFFFE5EAAAB7EEB6AAAAAAAAAAAAAAAAAAB36E7CEB0ABFFFFFFFFFFFF),
    .INIT_01(256'hEBE57EBFFFFE7EAAAF7EEB7AAAAAAAAAAAAAAAAAAB898F7EAD2BFFFFFFFFFFFF),
    .INIT_02(256'hEAFE1EBEFFFF7AAAADBFFAFAAAAAAAAAAAAAAAAAAACB3E3AABCFFFFFFFFFFFEF),
    .INIT_03(256'hFAFBEFEEFFF9BAAAACBBF9AAAAAAAAAAAAAAAAAAAAB2E8BAAAC6FFFFFFFFFE9A),
    .INIT_04(256'hAFFFBBBEFFEBBAAAACFBB8AAAAAAAAAAAAAAAAAAAAB8EFEAAAC0BFFFFFFFFFC2),
    .INIT_05(256'hDBFBEBBBFFF52AAAACFB6CEAAAAAAAAAAAAAAAAAAAACA3AAAAF46FFFFFFFFFA5),
    .INIT_06(256'hE7FBFAFFBF95EAAAACBB7BEAAAAAAAAAAAAAAAAAAAADEFAAAABC5BFFFFFFFFBA),
    .INIT_07(256'hFEF9FAEEBED7AAAAA8BF24EAAAAAAAAAAAAAAAAAAAAA6FAAFEAF1AFFFFFEBFFF),
    .INIT_08(256'hFDFF3EEFBFDBAAAAA8FF327AAAAAAAAAAAAAAAAAAAAA2AAEAEAB5FFFFFF97BFF),
    .INIT_09(256'hFF6F8BBFFE9EAAAAA8EF74AAAAAAAAAAAAAAAAAAAAAA3AA88BFB5EFFFFFD57BF),
    .INIT_0A(256'hFFFFA6FBFE2AAABFA9EE653AAAAAAAAAAAAAAAAAAAAA3AE27AAE86FFFFFF3C7A),
    .INIT_0B(256'hFFDFE6BBBFFAAA0EB9ED9F1FAAAAAAAAAAAAAAAAAAAAAB99EAAAC1BFFFFACBC3),
    .INIT_0C(256'hFFE3F5AFF93AAAAF02E88A86EAAAAAAAAAAAAAAAAAAAAD67AAAAB4AFFFFFF2FD),
    .INIT_0D(256'hFFFAE57AF93AAFFFA2EC8EF5EAAAAAAAAAAAAAAAAAAAB55EAAAAB0EFFFFFECBF),
    .INIT_0E(256'hFFFCBD9EF9EAB3ABFDA85EB5FAAAAAAAAAAAAAAAAAAAC97AAAAAB0FFFFFFFF2F),
    .INIT_0F(256'hFFFF7B7FFCAAC00042A442F97AAAAAAAAAAAAAAAAAAA35EAAAAAA86FFFFFFEDF),
    .INIT_10(256'hFFFF3B9ABCEAC09442E57C7D5EAAAAAAAAAAAAAAAAA89AAAAAAAAC3BFFFFFFA3),
    .INIT_11(256'hFFFF8FA46CEAC2BEF1E47ECF5BAAAAAAAAAAAAAAAAE66EAAAAAAAA7BFFFFFFE8),
    .INIT_12(256'hFFFFEAF25CEAC3FFE9F547E067AAAAAAAAAAAAAAAB89EAAAAAAAAA7BFFFFFFF8),
    .INIT_13(256'hFFFFF6EF98EAD3FFF9E001FF59EAAAAAAAAAAAAAAF27AAAAAAAAAA0BFFFFFFFE),
    .INIT_14(256'hFFFFFA96F5EAD7FFF9A5F41BC5BAAAAAAAAAAAAAB48AAAAAAAAAAB1FFFFFFFFF),
    .INIT_15(256'hFFFFFED4F0EAD3FFF994FA40F33AA8AAAAAAAAAAD63EBFFFAAAAAA9FFFFFFFFF),
    .INIT_16(256'hFFFFFF99E9EAD7FFFD99FF942D9EA8EAAAAAAAAB6955540FAAFAAA9BFFFFFFFF),
    .INIT_17(256'hFFFFFF99ECAAD7FFFCCEFFF90EDBAFEAAAAAAAACA40FAAAAABFAAA8BEEAFFFFF),
    .INIT_18(256'hFFFFFFD83DAADBFFFE8FFFEF9463A6AAA2AAAAE25FFABEAFFE9AAACF6FBFFFFF),
    .INIT_19(256'hFFFFFFFF6DFADBFFFF5FFE2BFD39E2AAF7AAAB8E610000001BEAAACA61EFFFFF),
    .INIT_1A(256'hFFFFFFDF1F7ACBFFFE2FFEBEFD0CA3AACAAAAE3140041404017EAADA4D2FFFFF),
    .INIT_1B(256'hFFFFFFFE5E3ACBFFFF7FFDFBFE0F23AA8AAAA990006FFFFF941BAAD62E7FFFFF),
    .INIT_1C(256'hFFFFFFECC33AC7FFFF7FF9FEFF074FAA8EAAFB44BAABFFFFEE03AAD97B3FFFFF),
    .INIT_1D(256'hFFFFFFEAF77AD3FFFF2FFBBEFFD5CBAACEAB782AAFFFFFFEBF0BAA9DA92BFFFF),
    .INIT_1E(256'hFFFFFFE8B53AF3FFFF7FFBBBFFD49FAADEB9D2BD9BFFFFFFFC1EAA9DB16BFFFF),
    .INIT_1F(256'hFFFFFFD8BC2AA7FFFFBFF9ABFFC11BAB5EE71AF9FBFFFFFFF83EAAFDE7EBFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_008192_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n653,addra[14:13]}),
    .dia({open_n657,open_n658,open_n659,open_n660,open_n661,open_n662,open_n663,1'b0,open_n664}),
    .rsta(rsta),
    .doa({open_n679,open_n680,open_n681,open_n682,open_n683,open_n684,open_n685,open_n686,inst_doa_i1_002}));
  // address_offset=8192;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h77CDD5F4A003628AAB579C4AAAAAAAAAAAAAAAAAAA5882128548080000000000),
    .INIT_01(256'hF77E05760803D2AAABD79C6AAAAAAAAAAAAAAAAAA83ABE7AA35C0A0000000000),
    .INIT_02(256'h55F7F77F8800E2AAAB14264AAAAAAAAAAAAAAAAAAA10724AA870000000000038),
    .INIT_03(256'h15F775BD880F2AAAA31E0D2AAAAAAAAAAAAAAAAAAA8629AAAA1F00000000019A),
    .INIT_04(256'hBFFF7FCF8AB31AAAA1942DA2AAAAAAAAAAAAAAAAAAA9072AAA3BC0000000003A),
    .INIT_05(256'hF7F77FC528076AAAA3BC6922AAAAAAAAAAAAAAAA2A8B86AAA2837000000000D5),
    .INIT_06(256'hDD70FD6168F8AAAAABF6E9AAAAAAAAAAAAAAAAAAAAA1662AAA25DC000000004C),
    .INIT_07(256'hFA75B5F9E91AAAAA81D8572AAAAAAAAAAAAAAAAAAAAAEEA2A2215B000283C800),
    .INIT_08(256'hFD3CCDD8CA32AAAAA15244CAAAAAAAAAAAAAAAAAAAAA6228AE88F8000000CC80),
    .INIT_09(256'hFDDD37528912AAAAA170692AAAAAAAAAAAAAAAAAAAAA4A8119D8C300000016C0),
    .INIT_0A(256'hFF9545F6A162A082ABD2C572AAAAAAAAAAAAAAAAAAA8E0AEEA84230000A243C5),
    .INIT_0B(256'hFFF1C4F6E2CA0A548BF93EFE2AAAAAAAAAAAAAAAAAA800398A283340000717B6),
    .INIT_0C(256'hFFD7E7BCAD4A82255CFD909EA8AAAAAAAAAAAAAAAAA0A94EAAAA83B0000A0FF2),
    .INIT_0D(256'hFFF057CD8E6A88002C3BB21FAAAAAAAAAAAAAAAAAAAAA75AAAAAA790000A33FD),
    .INIT_0E(256'hFFF7DB318FCA37A80511F80D48AAAAAAAAAAAAAAAAA0934AAAAA8608000A087F),
    .INIT_0F(256'hFFFE7E4289AA100A3497DC2BCAAAAAAAAAAAAAAAAAA8F5AAAAA88278000A8317),
    .INIT_10(256'hFFFF46BFCBAAB1B5A03DE743DAAAAAAAAAAAAAAAAA89B8AAAAA8A38E0000AAEF),
    .INIT_11(256'hFFFFFEE5730A326B8531EAF6D0AAAAAAAAAAAAAA2A284AAAAAAAAAA400008A33),
    .INIT_12(256'hFFFFC926390A30801123AE8FE4AAAAAAAAAAAAAA2891AAAAAAAAAA8400000084),
    .INIT_13(256'hFFFFF58C212A03DFF5AD406B2B2AAAAAAAAAAAAAA164AAAAAAAAA89400000001),
    .INIT_14(256'hFFFFF4D6BB2A0BFFF6C60000B70AAA2AAAAAAAAA87300AAAAAAAA84000000000),
    .INIT_15(256'hFFFFFE370D2227FFFC5D7C03AECAABAAAAAAAAAA1EC2AAAAAAAAA8B88000000A),
    .INIT_16(256'hFFFFFD18008227FFF659FFF08192A12AAAAAAAA8C0602BDD220AA89C22800000),
    .INIT_17(256'hFFFFFFC2C3280FFFF59AFFFDAE3A8D2AA2AAA0A9A1FFA0A2A17AAA1411F00000),
    .INIT_18(256'hFFFFFFF1410803FFFEB7FF7779F4862AA4AAA82C72009682A292AA30F8600000),
    .INIT_19(256'hFFFFFFF729CA0BFFFE5FFFC3D2A12EAA1CAAA8B0E42000025A8AAA125E100000),
    .INIT_1A(256'hFFFFFFDDD34A3BFFFDCFFE19FD97AEAABA2AA06C8009D75A0268A21ADDFA0000),
    .INIT_1B(256'hFFFFFFD5404233FFFD0FFD36FD20C4AA10AA89E00942AAAA9802AA3428000000),
    .INIT_1C(256'hFFFFFFED566A1FFFFDAFFD9C7F41D4AA1AAA1A09AD76A0081A04AA1B68600000),
    .INIT_1D(256'hFFFFFFE17B4ABFFFFFFFFD1EFF0BC2A8F2826A67FFFFF55F4A82AA3B0BE40000),
    .INIT_1E(256'hFFFFFFC174EAB7FFFF5FF7A5FF6E74A872A99E55BFFFFFFFFA00AA39AD640000),
    .INIT_1F(256'hFFFFFFF177A2A3FFFFDFF7897FF5F0A8F2A67D7B73FFFFFFFF12AAB9AA440000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_008192_003 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n712,addra[14:13]}),
    .dia({open_n716,open_n717,open_n718,open_n719,open_n720,open_n721,open_n722,1'b0,open_n723}),
    .rsta(rsta),
    .doa({open_n738,open_n739,open_n740,open_n741,open_n742,open_n743,open_n744,open_n745,inst_doa_i1_003}));
  // address_offset=8192;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h5D2915575FFF8FDFFCB5573FFFFFFFFFFFFFFFFFFF2953EFD057F7FFFFFFFFFF),
    .INIT_01(256'h55D23F57F7FF27FFFEB75D3FFFFFFFFFFFFFFFFFFDECE98FF49FF5FFFFFFFFFF),
    .INIT_02(256'hD55D8F5577FD3FFFFCF7FD9FFFFFFFFFFFFFFFFFFF47071FFDAFFFFFFFFFFFFF),
    .INIT_03(256'hF555F5F777FCFFFFF67DFEFFFFFFFFFFFFFFFFFFFFF17C7FFFCBFFFFFFFFFFC5),
    .INIT_04(256'h55555577757CEFFFF67FFCFFFFFFFFFFFFFFFFFFFFF4527FFF40FFFFFFFFFFC9),
    .INIT_05(256'h655D55FDD7FABFFFF4D7967FFFFFFFFFFFFFFFFFFFFE73FFF7D83FFFFFFFFFD8),
    .INIT_06(256'hFB57557D57C2FFFFFE57B67FFFFFFFFFFFFFFFFFFFF633FFFFF2AFFFFFFFFFFF),
    .INIT_07(256'hF5DCD5555741FFFFDEDFB27FFFFFFFFFFFFFFFFFFFFD33FFF7F627FFFD7FF7FF),
    .INIT_08(256'hFED59577F5EFFFFFF65DB19FFFFFFFFFFFFFFFFFFFFF177DF1DDA7FFFFFEBF7F),
    .INIT_09(256'hFD17ED5D77C7FFFFFCFD1257FFFFFFFFFFFFFFFFFFFF9FD44E2D07FFFFFE09FF),
    .INIT_0A(256'hFFCDDB555F37FFD7F4FD108FFFFFFFFFFFFFFFFFFFFD3FD33FDB4BFFFF5D3617),
    .INIT_0B(256'hFFEF79DD5F1FFF2356DE61A9FFFFFFFFFFFFFFFFFFFFFD4CDFFF607FFFFF4F6B),
    .INIT_0C(256'hFFD152F75E1FFFD88BDE6D4BFFFFFFFFFFFFFFFFFFFFF6B3FFFFF27FFFF5D1F6),
    .INIT_0D(256'hFFFFDA9D7E9FD5557BD6476AFFFFFFFFFFFFFFFFFFFFF20FFFFFF8FFFFF5F47F),
    .INIT_0E(256'hFFFEDCED7C1F6277707CA5F89DFFFFFFFFFFFFFFFFF5C61FFFFFD0F7FFF5FDBF),
    .INIT_0F(256'hFFFDB5BD7C7F600281FA037E9FFFFFFFFFFFFFFFFFFF88FFFFFFD4B7FFF57F47),
    .INIT_10(256'hFFFF17EFF6FFE06001D2BAB40FFFFFFFFFFFFFFFFFD665FFFFFFF6B5FFFF55F9),
    .INIT_11(256'hFFFF67F8B65F617FF2D2178385FFFFFFFFFFFFFFFF7B17FFFFFFFF1FFFFF75F6),
    .INIT_12(256'hFFFFFFF9A45F61FFDEF8A3789BFFFFFFFFFFFFFFFD647FFFFFFFFFBFFFFFFF75),
    .INIT_13(256'hFFFFF9DBC67F69FFF6FAA2148E7FFFFFFFFFFFFFF43BFFFFFFFFFF27FFFFFFFD),
    .INIT_14(256'hFFFFFD696A7F63FFFE5AD00FCADFFDFFFFFFFFFFD84D5FFFFFFFFD8FFFFFFFFF),
    .INIT_15(256'hFFFFFF605A7F43FFFEEAD500D93FFEFFFFFFFFFF4B17FFFFFFFFFD677FFFFFF5),
    .INIT_16(256'hFFFFFF6ED6FF43FFF646FD601CC7F67FFFFFFFFDBC0808AA5F5FFDEFDD7FFFFF),
    .INIT_17(256'hFFFFFF44947F6BFFFE67FFF683CFD07FFFFFFFFED288DFFD560FFFCDFF5FFFFF),
    .INIT_18(256'hFFFFFFE694DF67FFFF65FFFF6211DB7FD9FFFF512577415F574FFF473FDFFFFF),
    .INIT_19(256'hFFFFFFC2969F67FFFF8FFD1FDE3E79FF49FFFDED1AA000088F5FFF6D187FFFFF),
    .INIT_1A(256'hFFFFFFC8AC9F67FFFF9FFD75F60E5BFFEFFFF73A0008828002BFFF4D0835FFFF),
    .INIT_1B(256'hFFFFFFC88D1F47FFFD9FFE77FF8511FFEFFFD46008BFFFFD4027FF49153FFFFF),
    .INIT_1C(256'hFFFFFFD023BF6BFFFF3FF6FFFFA381FF6FFF4F02D7D7FFF7DF81FF641DBFFFFF),
    .INIT_1D(256'hFFFFFFFC223FC3FFFF3FFE5D7F6A4FFD27D79EB5FFFFFFF77D27FF4ED61FFFFF),
    .INIT_1E(256'hFFFFFFFC2A1FCBFFFF1FFC547F40C9FD07D4435EC7FFFFFFDF27FF44DA1FFFFF),
    .INIT_1F(256'hFFFFFFEC2097D1FFFF7FFC7CFFE22DFD87F30FF477FFFFFFFC07FFC45B9FFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_008192_004 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n771,addra[14:13]}),
    .dia({open_n775,open_n776,open_n777,open_n778,open_n779,open_n780,open_n781,1'b0,open_n782}),
    .rsta(rsta),
    .doa({open_n797,open_n798,open_n799,open_n800,open_n801,open_n802,open_n803,open_n804,inst_doa_i1_004}));
  // address_offset=8192;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hA9AEBFBEFFFFB12552AC97155555555555555555501C87606746FFFFFFFFFFFF),
    .INIT_01(256'hFA9E79FEFAFE895551EE8F15555555555555555556AD06755D4FFBFFFFFFFFFF),
    .INIT_02(256'hBFEC2D6CBEFE8555552AEC355555555555555555549D6B21571BBFFFFFFFFFAF),
    .INIT_03(256'hBFFE9EDCABEFC5555AB7BED55555555555555555555CD0015533BFFFFFFFFFB0),
    .INIT_04(256'h5FFEFE68BFE0A1555BE71E5555555555555555555558FC9555A0BFFFFFFFFFD4),
    .INIT_05(256'hEEF3FB67BFAED5555EB38AD55555555555555555555340555D0DBFFFFFFFFF8B),
    .INIT_06(256'hDFEFBFEE6FA845554023509155555555555555555559B9555558ABFFFFEFFEFD),
    .INIT_07(256'hB9B3BB896EE51555717A2D955555555555555555555279500C48A7FFFFBEEFFE),
    .INIT_08(256'hBEFC0FCFAFBD555154AE24A55555555555555555555200C4FC22BFFFFFE7FBBF),
    .INIT_09(256'hFFBB56FBAF0D55514ACFFC2C55555555555555555552A5769EF70FFFFFFA3EFF),
    .INIT_0A(256'hFF8B19A6FFE9553C4B88C105555555555555555555501528044C2BFFFFFB2DF7),
    .INIT_0B(256'hFEFE9936BC25520E7B9B5B631555555555555555555542E02500B37FFFFEC791),
    .INIT_0C(256'hFFEAAF1AFAA5511A50DC573B1555555555555555555549915555563FFFFFF1EE),
    .INIT_0D(256'hFFF1EFE4AEE53AFF98DE6C8E1555555555555555555503455555412FFFFFFC3E),
    .INIT_0E(256'hFFF96E6CFEA5C4B5BD40AE086355555555555555554A666555556DBFFFFFFE1F),
    .INIT_0F(256'hFFFEE2BFFB159000B949A18AC05555555555555555404815555564AFFFFFFFFB),
    .INIT_10(256'hFFFF8A7AB9050038D08E8A4C455555555555555555753B5555555D2BFFFFFFC3),
    .INIT_11(256'hFFFF4AEFF8E5916FBE84897CCA5555555555555555A40C55555556FBFFFFFFE5),
    .INIT_12(256'hFFFFC5811EE582FFC2AF40DF8815555555555555529C5155555554CAFFFFFEF5),
    .INIT_13(256'hFFFFAD93778596BAA29113BF67C55555555555555E990555555555D2FFFFFFFC),
    .INIT_14(256'hAABFF074DA958FFFF35EF40E2AB154155555555437A2B455555556EFFFFFFFFF),
    .INIT_15(256'hFFFFFDB6E59597FFF32DA0C26FD555155555555588AC5455055157BFFFFFFFFE),
    .INIT_16(256'hFFFFFE2374119FFFFE63FF78940950C555555547C474028215F557BBBFFFFFFF),
    .INIT_17(256'hFFFFFF556B159BFFF89DFBF200BD2FD5555555175392D55447B5557BAFFFFFFF),
    .INIT_18(256'hFFFFFFF32DF587FFFD0EFB7A7C9E3695435554CB6B97FAD0A87155A8FBFFFFFF),
    .INIT_19(256'hFFFFFEC0CD2597FFFFFFFD53EB248955F715538D3C8000061CF555B587BFFFFF),
    .INIT_1A(256'hFFFFFFCE1B2593FFFD0FFFF8FE490C556C155FB2C0152959034555C8B53FFFFF),
    .INIT_1B(256'hFFFFFFCE7525B7FFFFBFF438FD1C825535553C70119ABFFB6C3855CCFD6FFFFF),
    .INIT_1C(256'hFFFFFFCFED91EBFFFFAFF1FCBF4FAE542555A788A517AFEED80B45C3261BFFFF),
    .INIT_1D(256'hFFFFFFDA84005BFFFF4FF8FDFFFAFD56B97860158FFFEFE87B405583618BFFFF),
    .INIT_1E(256'hFFFFFFCF908527FFFFFFFC42BFF32F568831E161A3FFFFFFFB1D55DD6D5BFFFF),
    .INIT_1F(256'hFFFFFFFB8C9916FFFF2FF942BFC4FF5718122DBCD7FFFFFFF42D544CBC0FFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_008192_005 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n830,addra[14:13]}),
    .dia({open_n834,open_n835,open_n836,open_n837,open_n838,open_n839,open_n840,1'b0,open_n841}),
    .rsta(rsta),
    .doa({open_n856,open_n857,open_n858,open_n859,open_n860,open_n861,open_n862,open_n863,inst_doa_i1_005}));
  // address_offset=8192;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hBBCEEBE900018FAAACEB2C6AAAAAAAAAAAAAAAAAAB46FDFBA7D1000000000000),
    .INIT_01(256'hABB9DAE80500CAAAADE8213AAAAAAAAAAAAAAAAAAB22731EA8B4040000000000),
    .INIT_02(256'hAABBFBBB0101EAAAAD29143AAAAAAAAAAAAAAAAAAA974D2EAA25400000000045),
    .INIT_03(256'h3AABBB7E14162AAAAB2C477AAAAAAAAAAAAAAAAAAAAEBCFEAAE94000000001A1),
    .INIT_04(256'h2EABABDF00000EAAAB6857AAAAAAAAAAAAAAAAAAAAB1B0AAAAB6000000000034),
    .INIT_05(256'hFFAAAACE405FAAAAAF7DC6EAAAAAAAAAAAAAAAAAAAABE3AAAAE7C0000000006A),
    .INIT_06(256'hFBB0EA928026FAAAAFF984AEAAAAAAAAAAAAAAAAAAA953AAAAB3F00000100004),
    .INIT_07(256'hF4AA7AF2C16AEAAAAAE5DBAAAAAAAAAAAAAAAAAAAAAD17ABFFA8B10000001001),
    .INIT_08(256'hFE3EEEB01067AAAAAFA0D8AAAAAAAAAAAAAAAAAAAAAC6BAF07FAE4000010C000),
    .INIT_09(256'hFEFF3FA4110AAAAAB3F0921EAAAAAAAAAAAAAAAAAAACEABB141F31000005A800),
    .INIT_0A(256'hFF4A8AF801CEAAFFB2E4808AAAAAAAAAAAAAAAAAAAAE7A983FA694000005C3D9),
    .INIT_0B(256'hFFF2C8F8402AAD01F6F632B6AAAAAAAAAAAAAAAAAAAAAA71FABEB38000012B3D),
    .INIT_0C(256'hFFEB8B7D02AAAAA508F73AB8EAAAAAAAAAAAAAAAAAAAA9D7AAAAAC1000004FF1),
    .INIT_0D(256'hFFF0ABCF15EABAFFEC346A8EAAAAAAAAAAAAAAAAAAAAE24EAAAABF10000013FE),
    .INIT_0E(256'hFFFBF733073AC41EB522EFBD2AAAAAAAAAAAAAAAAAABF36AAAAAA940000004BF),
    .INIT_0F(256'hFFFCBD8007EAA0007C6BE7B2EEAAAAAAAAAAAAAAAAAFC9AAAAAAB8800000012F),
    .INIT_10(256'hFFFFA97006EAA36B013BA37D4AAAAAAAAAAAAAAAAABF63AAAAAAAB540000005F),
    .INIT_11(256'hFFFFF96F82EAB1955E3EEF2692AAAAAAAAAAAAAAAA8C7EAAAAAAAC1400000002),
    .INIT_12(256'hFFFFC60FF7EAB040221346FF9FEAAAAAAAAAAAAAAA75BAAAAAAAAB1400000109),
    .INIT_13(256'hFFFFFA4782AAA3EFFA5EC06C96AAAAAAAAAAAAAAA9DEFAAAAAAAAA6800000002),
    .INIT_14(256'hFFFFF8F787AAA7FFF9C90C36BB7AABAAAAAAAAAAA66FAAAAAAAAAAC000000000),
    .INIT_15(256'hFFFFFD33AEAABBFFFCAEBC03ECFAA8EAAAAAAAAA89BBABFFFAAAAB2400000000),
    .INIT_16(256'hFFFFFE31BAEEBBFFF9A6FEE03D4EA8EAAAAAAAABD73ABA80AEFAAA3040000000),
    .INIT_17(256'hFFFFFFFB2AAABFFFFA65FFFB5023B4EAAEAAAAAE4F903AAFAD1AAAA510000000),
    .INIT_18(256'hFFFFFFEAFD3AA3FFFD7BFF9FA3EAB1EAB3AAAAED7BFD142EFB9AAAB5C4400000),
    .INIT_19(256'hFFFFFFCC2D2AA7FFFDAFFE97E015BBAAC7AAAB345A000004C2BAAAA0A9500000),
    .INIT_1A(256'hFFFFFFD18D6AB7FFFECFFEF7FE2BAFAAE7AAADDC0006EBA5016EAAC8F4800000),
    .INIT_1B(256'hFFFFFFC07E6AA3FFFE0FFF39FF02F6AAAAAAB1D0028155556413AAD94BD00000),
    .INIT_1C(256'hFFFFFFD13BFAEFFFFE5FFFF8FFC2A2ABBEAA85069AB95004354AAAD32AC40000),
    .INIT_1D(256'hFFFFFFC4183ACBFFFFFFF6EDFF52D3AB2AAF448B7FFFFAAF905FAA96E9940000),
    .INIT_1E(256'hFFFFFFC507EACBFFFFAFF29EBF81B3AB0ABC69ABBFFFFFFFE72AAAD0AC440000),
    .INIT_1F(256'hFFFFFFE1003EFBFFFFEFF3EEFFE4A3AB4B95B6FAA7FFFFFFFF1EAAC0C7040000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_008192_006 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n889,addra[14:13]}),
    .dia({open_n893,open_n894,open_n895,open_n896,open_n897,open_n898,open_n899,1'b0,open_n900}),
    .rsta(rsta),
    .doa({open_n915,open_n916,open_n917,open_n918,open_n919,open_n920,open_n921,open_n922,inst_doa_i1_006}));
  // address_offset=8192;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hAE162BABFFFF4FFFFF3AEBFFFFFFFFFFFFFFFFFFFFA2A2DFE9AFFFFFFFFFFFFF),
    .INIT_01(256'hAAE16FEAFFFE2BFFFE7AEAFFFFFFFFFFFFFFFFFFFFC98AEFFB6FFFFFFFFFFFFF),
    .INIT_02(256'hEAAE4FAAFFFE2FFFFFFBFFBFFFFFFFFFFFFFFFFFFFABBBAFFE9FFFFFFFFFFFEF),
    .INIT_03(256'hEAAAFAFBFFFCAFFFF8BFFCFFFFFFFFFFFFFFFFFFFFF3BEBFFFD3FFFFFFFFFF0E),
    .INIT_04(256'hAAAAAABBFFEEBFFFF9BFFDFFFFFFFFFFFFFFFFFFFFFEBABFFF91BFFFFFFFFFC7),
    .INIT_05(256'h9EAEAAFAFFF07FFFFDEB78FFFFFFFFFFFFFFFFFFFFF9BBFFFFF02FFFFFFFFFE4),
    .INIT_06(256'hE6ABAABEBF90FFFFFCAB2ABFFFFFFFFFFFFFFFFFFFFBBBFFFFFC5BFFFFFFFFFF),
    .INIT_07(256'hFAECEAAEBF83FFFFFCEF70BFFFFFFFFFFFFFFFFFFFFFFBFFFFFA1FFFFFFEBFFF),
    .INIT_08(256'hFDEA6ABFBFDFFFFFF8AF726FFFFFFFFFFFFFFFFFFFFEBBFEAAFE1BFFFFFD7BFF),
    .INIT_09(256'hFE3ADAAFFFFBFFFFF9BE21BFFFFFFFFFFFFFFFFFFFFE6FF9EFABDBFFFFFD07BF),
    .INIT_0A(256'hFFEEE7ABFF6FFFFFFCFF6F6FFFFFFFFFFFFFFFFFFFFEBFB3FFEB96FFFFFE392B),
    .INIT_0B(256'hFFDFB6EFFEAFFFBBBDED9E5AFFFFFFFFFFFFFFFFFFFFFE8FFFFF80BFFFFF8FD7),
    .INIT_0C(256'hFFE2F1FBF96FFFEEE7EDCFD6FFFFFFFFFFFFFFFFFFFFFB2FFFFFF4FFFFFFE2F9),
    .INIT_0D(256'hFFFFE56EFD6FFAFFF3E88BA1BFFFFFFFFFFFFFFFFFFFEDFFFFFFF0BFFFFFF8BF),
    .INIT_0E(256'hFFFDECDEFCFFEAFBABBC5BF3AFFFFFFFFFFFFFFFFFFFD9AFFFFFE4FFFFFFFE7F),
    .INIT_0F(256'hFFFF7A7FFDBF800116F51AB93FFFFFFFFFFFFFFFFFFF27BFFFFFF86FFFFFFF8B),
    .INIT_10(256'hFFFF2BDAB9FF909002E06DFBFBFFFFFFFFFFFFFFFFF89FFFFFFFF87FFFFFFFF6),
    .INIT_11(256'hFFFF9FC169FF82BFE5E53B9A7EFFFFFFFFFFFFFFFFA3EFFFFFFFFE2FFFFFFFE9),
    .INIT_12(256'hFFFFFFE219FF82FFEDF45EA563FFFFFFFFFFFFFFFECFFFFFFFFFFF7FFFFFFFFB),
    .INIT_13(256'hFFFFF6EAC8BF86FFF9F550AB0DBFFFFFFFFFFFFFFA73FFFFFFFFFF5BFFFFFFFE),
    .INIT_14(256'hFFFFFE8EA4BF83FFFDA5E41F95FFFEFFFFFFFFFFECCFFFFFFFFFFE4FFFFFFFFF),
    .INIT_15(256'hFFFFFF8DA0BF93FFFDD5EA01F27FFFFFFFFFFFFFB72BFFFFFFFFFFDBFFFFFFFF),
    .INIT_16(256'hFFFFFF8CF8FF93FFF989FF902FFBFBFFFFFFFFFF29C5513BABFFFF8BFFFFFFFF),
    .INIT_17(256'hFFFFFF98A9BF97FFFD9BFFFD4BCBFAFFFBFFFFFCE52BAFFAAEAFFFDEFFFFFFFF),
    .INIT_18(256'hFFFFFFD92EFF8BFFFF9AFFAF9026FFFFEFFFFFF7CEBBEBEEABBFFF9B2FFFFFFF),
    .INIT_19(256'hFFFFFFEE7FAF8BFFFF4FFF3FED7BB2FFEFFFFF8AF01000003ABFFF8F24BFFFFF),
    .INIT_1A(256'hFFFFFFFE7AEF8BFFFF6FFC3AF90CF7FFCFFFFF750004414000EFFFF31B6FFFFF),
    .INIT_1B(256'hFFFFFFEEDEAF9BFFFE6FF9FAFE4A6AFFDFFFFF90007FFFFE800FFFF67A7FFFFF),
    .INIT_1C(256'hFFFFFFEF977FC7FFFF3FFD3EFF135AFF9FFFAB012BEBFFFBFF46FFFCEE2FFFFF),
    .INIT_1D(256'hFFFFFFFEA6FFF3FFFF3FF87FBFC59FFFCBFFEC7BBFFFFFFBAE0BFFBDBF3FFFFF),
    .INIT_1E(256'hFFFFFFFFAD7FF3FFFF2FF87CFF8DCFFFBBFB97A85BFFFFFFED0BFFFBE3FFFFFF),
    .INIT_1F(256'hFFFFFFDBAB2FE6FFFFBFF950FFDF1FFFFBAF0FF1EBFFFFFFFC2FFFEBB3BFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_008192_007 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n948,addra[14:13]}),
    .dia({open_n952,open_n953,open_n954,open_n955,open_n956,open_n957,open_n958,1'b0,open_n959}),
    .rsta(rsta),
    .doa({open_n974,open_n975,open_n976,open_n977,open_n978,open_n979,open_n980,open_n981,inst_doa_i1_007}));
  // address_offset=16384;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFE0C81EA6EFFFFFF200FFD0C3EEF78D4FEEBFFFFFFFFE2BFAC6C01BFFFF),
    .INIT_01(256'hFFFFFFC9E946EBEFFFFFF609FFC813AA7ADA3FFFF3FFFFFFF40BFAD0734BFFFF),
    .INIT_02(256'hFFFFFFCCD162FCFFFFFFFE9BBFF94274BB26FFE8BBFFFFFFF43BFEA8CE3BFFFF),
    .INIT_03(256'hFFFFFFFC92A6F73FFFFFFF3EBFDDAE8DE197FFD126FFFFFFF3EBFE367E3BFFFF),
    .INIT_04(256'hFFFFFFF265A6BF4FFFFFFFFFFFFF6DF29D7FFFF007FFFFFFE63BFF6D36E2AFFF),
    .INIT_05(256'hFFFFFFF7254FBBA3FFFFFFFFFE7A7BE0F663FFE01BFFFFFFF7AFFF152FF06BAA),
    .INIT_06(256'hFFFFFFFE5B9BAAECFFFFFFFFF9FABEFEE4DFFFD437FFFFFFDCABFE350CCA06F0),
    .INIT_07(256'hFFFFFFFF0CBBAABEBFFFFFFF97FAFFFAB2FFFFE47BFFFFFF2BAFEC48550B9AC0),
    .INIT_08(256'hFFFFFFFF1442AAAEB7FFFFFE5FFFFFFEBF9FEFFB5FFFFFFF5AAEE23779778BFF),
    .INIT_09(256'hFFFFFFFF4FDDAAAB862FFF0CEEFFFFFEFE9FFFFC7FFFFFFEFEAFEB5779CBCBFF),
    .INIT_0A(256'hFFFFFFFFF3D9AAAAB94D3B0BAABFFBFEBECFFFFFFFFFFFFF7EAFBAA08977F9BF),
    .INIT_0B(256'hFFFFFFFFE149AAAAAAA41EEAAABFFEFEBEE6FFFFFFFFFFFEBFEBA031DB2A29BF),
    .INIT_0C(256'hFFFFFFFFFD76AAAFFFFFFEABFABFFFBEBEBBFFFFFFFFFFF03FFBAF20D7476E7F),
    .INIT_0D(256'hFFFFFFFFFFE3FFFFFFFFFEBFFFFFFBFBFFFEBFFFFFFFFFD3FFFEFFB2BBA3EE7F),
    .INIT_0E(256'hFFFFFFFFFF08FFFFFFFFFFFFFFFFE5EBFFFB8BFFFFFFFFF6FFFA3A2331FA8B7F),
    .INIT_0F(256'hFFFFFFFFFF8DFFFFFFFFFFFFFFFF9DEBFFFAE7FFFFFFFF2EBFFBB61D44FB3AAE),
    .INIT_10(256'hFFFFFFFFFFB22FFFFFFFFFFFFFFF18AFFFFAB87FFFFFFD7EBFEA5B70F3FF6F6B),
    .INIT_11(256'hFFFFFFFFF2766FFFFFFFFFFFFFFF58BFFFFEEE07FFFFCEBBFFFD81038FFB1F4F),
    .INIT_12(256'hFFFFFFFF9F656BFFFFFFFFFAAAFB9DEBFFFFFB1C565CD6FBFFED0DC86FFFEFD1),
    .INIT_13(256'hFFFFFFFFC590EAFFFFFFFFFAAAFBD2FFFFFFFAEF44188BFFFFEDB351FFFFB3B3),
    .INIT_14(256'hFFFFFFCE07467AFFFFFFFFFFFFFFFBFEAAAAAAFEBEEBABFFFFE8BD6E3FFFE0EF),
    .INIT_15(256'hFFFFFF689F2A0ABFFFFFFFFAAAABFE082EBABABAAAAAABFFFFAA30A351ABFABE),
    .INIT_16(256'hFFFFFFFFFCD1DABFFFFFFFEABF0AE1F942B1E6FAFFFFFFFFFEABC6F540DAF93B),
    .INIT_17(256'hFFFFFFFFF8853ABFFFFFFF82C346C2965FF8207AFFFFEBFFFEFB3BFFFF6BAFDE),
    .INIT_18(256'hFFFFFFFF407BEEBFFFFFACE3C634AFFFFFFFF79EFFFFABFFFA9AB6FFFFE748EB),
    .INIT_19(256'hFFFFFFEFAD4F5ABFFFEE0389FFFFFFFFFFFFFF1BFFFFFFFFE9621CFFFFFE1A9B),
    .INIT_1A(256'hFFFFFE8E9DF7B2BFFFEAC3FFFFFFFFFFFFFFFF51EAFFFFFFEBB25CBFFFFFF8EE),
    .INIT_1B(256'h0550951A85D59FBFFFEAE3FFFFFFFFFFFFFFFF727AFFFFFFA2E983FFFFFFFFFF),
    .INIT_1C(256'h00C172955445F4AFFFAACAD8FFEC3BBA447CFF7B9AFFFFFFB7EA2CBFFFFFFFFF),
    .INIT_1D(256'hAAAA95554556ADEFFFE98F25555555D5555AA76636BFFFFEA17AB98FFFFFFFFF),
    .INIT_1E(256'h555555555556F5ABFEF8D9BFEAAAAAAAAABA9B6EBEAFFFFEACA8233EFFFFFFFF),
    .INIT_1F(256'h555555555552AC6BFEF82FFEAEAABBFFA16AEEBBC9AFFFEFD7C4730FFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_016384_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1007,addra[14:13]}),
    .dia({open_n1011,open_n1012,open_n1013,open_n1014,open_n1015,open_n1016,open_n1017,1'b0,open_n1018}),
    .rsta(rsta),
    .doa({open_n1033,open_n1034,open_n1035,open_n1036,open_n1037,open_n1038,open_n1039,open_n1040,inst_doa_i2_000}));
  // address_offset=16384;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFE0C9854DFFFFFFFB51FFDCB144AD91BBEDF2FFFFFFF84555471B415555),
    .INIT_01(256'hFFFFFFCCE89D4EFFFFFFFE5EFFF967247E54FFD9FAFFFFFFF8E55544C9415555),
    .INIT_02(256'hFFFFFFEDC0E956BFFFFFFDD7FFF007B641F8FFCDF6FFFFFFF455554A51315555),
    .INIT_03(256'hFFFFFFFD82695B7FFFFFFFAFFFE5971E62CBFFD0A3FFFFFFFD15550825315555),
    .INIT_04(256'hFFFFFFF622B955BFFFFFFFFFFF8414590927FFD143FFFFFFF685554435390555),
    .INIT_05(256'hFFFFFFFF6321557FFFFFFFFFFFD55540526FFFC153FFFFFFC155554C3528C500),
    .INIT_06(256'hFFFFFFFF1821555EFFFFFFFFFF555555517FFFF56BFFFFFFEE5555282230E3F1),
    .INIT_07(256'hFFFFFFFD9D3555563FFFFFFFF1555555517FFFE56FFFFFFFD15554283A317BBF),
    .INIT_08(256'hFFFFFFFFD1105554ABFFFFF855555555556FFFF6EFFFFFFF51545B030A691BFF),
    .INIT_09(256'hFFFFFFFFE5CA55550BBFFFD945555555557FFFFFFFFFFFFEC55552F3068168FF),
    .INIT_0A(256'hFFFFFFFFE24A555551AD5141555555555543FFFFFFFFFFFD45555660A2C957BF),
    .INIT_0B(256'hFFFFFFFFEF4E555554155155555555555559FFFFFFFFFFFB15554661819D90FF),
    .INIT_0C(256'hFFFFFFFFF0985555555555555555555555537FFFFFFFFFF195554CB08BEB04DF),
    .INIT_0D(256'hFFFFFFFFFE4D555555555555555554555554DFFFFFFFFFEC555551F28540346F),
    .INIT_0E(256'hFFFFFFFFFC7C55555555555555555155555537FFFFFFFFF05555A3A34956FCA3),
    .INIT_0F(256'hFFFFFFFFFEF955555555555555554C55555548FFFFFFFF21555508CCB6537B1F),
    .INIT_10(256'hFFFFFFFFFE2695555555555555554C155555523FFFFFFC8555544337E955EECC),
    .INIT_11(256'hFFFFFFFFFE4E95555555555555550D15555554FBFFFFEF155556740FA5554FE6),
    .INIT_12(256'hFFFFFFFFDD8A95555555555555550955555555D36EE0E4555555DC3F85557FF9),
    .INIT_13(256'hFFFFFFFC834F5555555555555555515555555546AEAD61555556B5AA555507F5),
    .INIT_14(256'hFFFFFF90EDDA155555555555555555555555555415415555555496C8955542FE),
    .INIT_15(256'hFFFFFFF83E92655555555555555554A2855015555555555555551A88DB5557FF),
    .INIT_16(256'hFFFFFFFFFDF8E5555555555555A051BEBFBE98555555555555556BFE3D75503F),
    .INIT_17(256'hFFFFFFFFFB23C5555555552847AD6EC5BBFA6C95555555555555B7FFF6F105FF),
    .INIT_18(256'hFFFFFFFFDAAE9555555504B96F4FBFFFFFFFFAA55555555554644AFFFF93066B),
    .INIT_19(256'hFFFFFFF69DDA115555546BD6BFFFFFFFFFFFFF215555555556A89DFFFFFF9EEB),
    .INIT_1A(256'hFFFFF9F9A76E3D5555548BFFFFFFFFFFFFFFFFDE55555555554E63FFFFFFFE43),
    .INIT_1B(256'h5555FB6A8BBF61555554CBFFFFFFFFFFFFFFFFC2955555555ACC1A3FFFFFFFFF),
    .INIT_1C(256'h00C05EBFEEEE6655555486E0AABC45145147BFC4E5555555597080FFFFFFFFFF),
    .INIT_1D(256'hAAAABFFFEFFC4E555556D6C55555555555506F9C6955555543903A7FFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFD1C155556910000000000000015B4145555554E099DBFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFD539555568000140011550A8104801E55555557FEC52BFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_016384_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1066,addra[14:13]}),
    .dia({open_n1070,open_n1071,open_n1072,open_n1073,open_n1074,open_n1075,open_n1076,1'b0,open_n1077}),
    .rsta(rsta),
    .doa({open_n1092,open_n1093,open_n1094,open_n1095,open_n1096,open_n1097,open_n1098,open_n1099,inst_doa_i2_001}));
  // address_offset=16384;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFDB372AB7FFFFFFF9AAFFE65AAB5E6C2FF2FFFFFFFFFD3AAAA9C3EBFFFF),
    .INIT_01(256'hFFFFFFE7173AB5FFFFFFF9A6FFE7CCDBC5F5BFF6FBFFFFFFF83AAAAA52EBFFFF),
    .INIT_02(256'hFFFFFFE33F5EA8FFFFFFFF7FFFEFECCF9F03FFF6FFFFFFFFF8AAAAB0369BFFFF),
    .INIT_03(256'hFFFFFFF37D5EACBFFFFFFFFFFFEB68F39873FFEABBFFFFFFF0EAAAB1D29BFFFF),
    .INIT_04(256'hFFFFFFF9DC4EAA2FFFFFFFFFFFFAEBA2F3DBFFEAABFFFFFFF1EAAAF7C29BAFFF),
    .INIT_05(256'hFFFFFFF8DD8EAA8BFFFFFFFFFFEAEABAADDBFFFABFFFFFFFF2AAAAE7C29B3FAA),
    .INIT_06(256'hFFFFFFFDE5CEAAA2FFFFFFFFFFAAAAAAAFBFFFFE9BFFFFFFC3AAAA93C78A095A),
    .INIT_07(256'hFFFFFFFF30CAAAA9FFFFFFFFFAAAAAAAAAAFFFFEDFFFFFFF9EAAAA87D38BCFEA),
    .INIT_08(256'hFFFFFFFF3CBBAAAB5BFFFFFFFAAAAAAAAAAFFFFD2FFFFFFFFEABAD9CD7DBA7FF),
    .INIT_09(256'hFFFFFFFFC827AAAAE1BFFFA7BAAAAAAAAABFFFFEBFFFFFFF3AAAAD1CDB6BE7FF),
    .INIT_0A(256'hFFFFFFFFD927AAAAAF03AEEEAAAAAAAAAAAFFFFFFFFFFFFEFAAAA95F4F3BFCFF),
    .INIT_0B(256'hFFFFFFFFF3E3AAAAABEFFAAAAAAAAAAAAAA3FFFFFFFFFFFCEAAABC1E7E37BA7F),
    .INIT_0C(256'hFFFFFFFFFFE3AAAAAAAAAAAAAAAAAAAAAAACFFFFFFFFFFFBEAAAB10F7C21AE3F),
    .INIT_0D(256'hFFFFFFFFFDB2AAAAAAAAAAAAAAAAAAAAAAAB3FFFFFFFFFE3AAAAA54D69EBDE9F),
    .INIT_0E(256'hFFFFFFFFFFF2AAAAAAAAAAAAAAAAAFAAAAAACFFFFFFFFFCBAAAAD51CF2FDE79F),
    .INIT_0F(256'hFFFFFFFFFF37AAAAAAAAAAAAAAAAB3AAAAAAB3FFFFFFFF9EAAAAD133CEF9BDF3),
    .INIT_10(256'hFFFFFFFFFF59EAAAAAAAAAAAAAAAF3EAAAAAACBFFFFFFE3AAAABC4CF1BFF3F37),
    .INIT_11(256'hFFFFFFFFF9D1EAAAAAAAAAAAAAAAF3EAAAAAAB0BFFFFE0EAAAAB4FEC6FFFAF89),
    .INIT_12(256'hFFFFFFFFE7B0EAAAAAAAAAAAAAAAB3AAAAAAAAF4ABAE0FAAAAAB73B0AFFFDBF3),
    .INIT_13(256'hFFFFFFFF6868AAAAAAAAAAAAAAAABEAAAAAAAAB90403BEAAAAA84EC2FFFFBBF9),
    .INIT_14(256'hFFFFFFE50329AAAAAAAAAAAAAAAAAAAAAAAAAAABEABEAAAAAAAA7B57BFFFEAFD),
    .INIT_15(256'hFFFFFF96EF38FAAAAAAAAAAAAAAAABFFFAAFEAAAAAAAAAAAAAAAAC712BFFFDFF),
    .INIT_16(256'hFFFFFFFFFE3A3AAAAAAAAAAAAAFFAB4000406FAAAAAAAAAAAAAAB1FC82FFFABF),
    .INIT_17(256'hFFFFFFFFFCE83AAAAAAAAAFFAC05416BAFFE92EAAAAAAAAAAAAAC7FEBD1FAF3F),
    .INIT_18(256'hFFFFFFFFA1976AAAAAAAFA4141BEFFFFFFFFF97AAAAAAAAAAB8B93FFFFF9BEDF),
    .INIT_19(256'hFFFFFFFD762FBEAAAAABC06EFFFFFFFFFFFFFF8EAAAAAAAAAB1F26FFFFFFA547),
    .INIT_1A(256'hFFFFFF47E4FBCEAAAAAB2BFFFFFFFFFFFFFFFFB3AAAAAAAAAA7DECFFFFFFFEBF),
    .INIT_1B(256'hAAAA40AFE2EACEAAAAAB3BFFFFFFFFFFFFFFFFB9EAAAAAAAAD36A9FFFFFFFFFF),
    .INIT_1C(256'hAA6ABBEAABBADFAAAAAB6FEE5556BFBFAABEFFBD3AAAAAAAAD5E867FFFFFFFFF),
    .INIT_1D(256'hFFFFEAAABAAAF3AAAAAB05100000000000055BB11EAAAAAAB8BA946FFFFFFFFF),
    .INIT_1E(256'hAAAAAAAAAAABF2EAAAAB045555555555555547914BAAAAAAB0A2B31FFFFFFFFF),
    .INIT_1F(256'hAAAAAAAAAAABF4EAAAAB1555540011550001515543AAAAAABD60398FFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_016384_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1125,addra[14:13]}),
    .dia({open_n1129,open_n1130,open_n1131,open_n1132,open_n1133,open_n1134,open_n1135,1'b0,open_n1136}),
    .rsta(rsta),
    .doa({open_n1151,open_n1152,open_n1153,open_n1154,open_n1155,open_n1156,open_n1157,open_n1158,inst_doa_i2_002}));
  // address_offset=16384;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFB574080FFFFFFF702FFCA4888D86ADFFCF3FFFFFFF48AA82324EC0000),
    .INIT_01(256'hFFFFFFCD55D285FFFFFFF50DFFFF7FB875987FE47DFFFFFFF4CAA8808ECC0000),
    .INIT_02(256'hFFFFFFD7779AA9FFFFFFFC5BFFD9C7BE8AFCFFE4F3FFFFFFF80AA82BB836AAAA),
    .INIT_03(256'hFFFFFFD5D792A1BFFFFFFF7FFFD14394BBFFFFC079FFFFFFF6AAA82E589E2AAA),
    .INIT_04(256'hFFFFFFFB5F72A87FFFFFFFFFFFC8CB0E3DFBFFC22BFFFFFFF92AA84B721ED200),
    .INIT_05(256'hFFFFFFFDD63A2A1FFFFFFFFFFF0AEA808F7FFFE213FFFFFFEA8AA843583668FF),
    .INIT_06(256'hFFFFFFFFF69AAA8DFFFFFFFFFC2A28AAAD8FFFE4BFFFFFFFFCAAA8BFD23FD9F2),
    .INIT_07(256'hFFFFFFFE5C3AAA8B3FFFFFFF60AAAAAAA21FFFFC5FFFFFFF42AAA0BDC6BCB5D5),
    .INIT_08(256'hFFFFFFFF7E38AAAAD7FFFFFCDAAAAAAAAA3FFFFB7FFFFFFF70A8A305E67CE7FF),
    .INIT_09(256'hFFFFFFFFB0C4AAA2855FFFE5AAAAAAAAAA0D7FF57FFFFFFFCAA8A365404C36FF),
    .INIT_0A(256'hFFFFFFFFFB84AAA2ABD72AC8AAAAAAAAAAAB7FFFFFFFFFFE4A8A8BB5DAC4037F),
    .INIT_0B(256'hFFFFFFFFDECCAAAAA82F700AAAAAAAAAAAACFFFFFFFFFFFD2A8A8795DA6ECC7F),
    .INIT_0C(256'hFFFFFFFFF186AAA0AAA82AA8AAAAAAAAAA813FFFFFFFFFF32AAA8E5DF1FFB3EF),
    .INIT_0D(256'hFFFFFFFFFD26AAAAAAAAAAAAAAAAA2AAAAAA4D7FFFFFFFDEAAAA2A7D483293BF),
    .INIT_0E(256'hFFFFFFFFFEEEAAAAAAAAAAAAAAAA87AAAAAA3B7FFFFFFFF2AAAA11754E01D4F3),
    .INIT_0F(256'hFFFFFFFFFDEF2AAAAAAAAAAAAAAA3D2AAAAAA6FFFFFFFF9AAAAA24F537AFB70D),
    .INIT_10(256'hFFFFFFFFFF99AAAAAAAAAAAAAAAA752AAAAA833FFFFFFEEAAAA8E95CFEA8DFEE),
    .INIT_11(256'hFFFFFFFFF5452AAAAAAAAAAAAAAAF52AAAAAA8FFFFFFF7AAAAAA15417008AFFB),
    .INIT_12(256'hFFFFFFFF64C52AAAAAAAAAAAAAAAB72AAAAAAA31BDFA76AAAAA33525D80217C5),
    .INIT_13(256'hFFFFFFFECB050AAAAAAAAAAAAAAA9CAAAAAAAA8173D702AAAAA1D415000A43F2),
    .INIT_14(256'hFFFFFFE85EEF8AAAAAAAAAAAAAA022AAAAAAAAAA28802AAAAAA8F0844AA8B3FF),
    .INIT_15(256'hFFFFFFF43F44CAAAAAAAAAAAAAAAA00028882AAAAAAAAAAAAAAA03ECC6A8097D),
    .INIT_16(256'hFFFFFFFFFC6C42AAAAAAAAAA8008837FFFDDEA2AAAAA0AAAAAAA8DF114A00E3F),
    .INIT_17(256'hFFFFFFFFF519E2AAAAAAAA008F723562FDF5B42AAAAAAAAAAAA81BFF79F2DA6F),
    .INIT_18(256'hFFFFFFFFC7F5CAAAAAA8AA5C17215FFFFFFFF7EAAAAAAAAAAA320DFFFFEB2197),
    .INIT_19(256'hFFFFFFD94CC71AAAAAAA5761FFFFFFFFFFFFFF38AAAAAAAAAAF066FFFFFD6577),
    .INIT_1A(256'hFFFFFC5C5B1D92AAAAAA6FFFFFFFFFFFFFFFFF7EAAAAAAAAA809517FFFFFFD01),
    .INIT_1B(256'h0AA07F3DCD7F12AAAA8AE7FFFFFFFFFFFFFFFFCB2AAAAAAAA1E6EDBFFFFFFFFF),
    .INIT_1C(256'h00C2A57FFFFF1CAAAA82E1FA5F5C22608029FFE24AAAAAAAA233FAFFFFFFFFFF),
    .INIT_1D(256'h55557FFFDFFFA6AAAAA869E00AAAA0000AA01F4432AAAAAA896FF59FFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFCA6AAAA8AC2202AAAAAAA8028227882AAAAAAAFDA467FFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFF4AB2AAA8A40A20BD7EE287FDEA2CA84AAAAAAB55DE21FFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_016384_003 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1184,addra[14:13]}),
    .dia({open_n1188,open_n1189,open_n1190,open_n1191,open_n1192,open_n1193,open_n1194,1'b0,open_n1195}),
    .rsta(rsta),
    .doa({open_n1210,open_n1211,open_n1212,open_n1213,open_n1214,open_n1215,open_n1216,open_n1217,inst_doa_i2_003}));
  // address_offset=16384;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFC40037DBFFFFFFFCFFFFDBA7DDA5B637FB75FFFFFFFCBFFDD4C39FFFFF),
    .INIT_01(256'hFFFFFFD20007DAFFFFFFFCF1FFF0A8E52AC8FFD3FDFFFFFFFC1FFD7F0B1FFFFF),
    .INIT_02(256'hFFFFFFDA2087F67FFFFFFDAFFFFE12C3C7A9FFD17DFFFFFFFCDFFD7CABED5555),
    .INIT_03(256'hFFFFFFFA8207F6FFFFFFFFFFFFDC3EC16EABFFDF5FFFFFFFF8FFFDD223EDD555),
    .INIT_04(256'hFFFFFFFC0227FD3FFFFFFFFFFFFF3CF16A27FFDDFFFFFFFFD87FFD12036DFDFF),
    .INIT_05(256'hFFFFFFFE02CF7F6FFFFFFFFFFF7FBFDDF00FFFDDEFFFFFFFD9DFFFB82147B7FF),
    .INIT_06(256'hFFFFFFFE8A67FFDBFFFFFFFFFDFFFFFFF2FFFFDBCFFFFFFFC9FFFD40096F06A5),
    .INIT_07(256'hFFFFFFFF20CFFFD6FFFFFFFFDFFFFFFFF7FFFFF9A7FFFFFFCFFFF54021EF677F),
    .INIT_08(256'hFFFFFFFF28E5FFFF0FFFFFF707FFFFFFFFDFFFFC3FFFFFFF25FFF440090FD3FF),
    .INIT_09(256'hFFFFFFFF66B9FFF7F87FFFF07FFFFFFFFFDFFFFDFFFFFFFD3FFFFE20251FF1FF),
    .INIT_0A(256'hFFFFFFFFEEB1FFF7FC085FBDFFFFFFFFFFDFFFFFFFFFFFFD1FFFDC80AF17FE7F),
    .INIT_0B(256'hFFFFFFFFDB39FFFFFD58075FFFFFFFFFFFD1FFFFFFFFFFF6FFFFD8A08F91FDBF),
    .INIT_0C(256'hFFFFFFFFFE7BFFFFFFFD7FFFFFFFFFFFFFDE7FFFFFFFFFFE7FFFD08086B27FBF),
    .INIT_0D(256'hFFFFFFFFFCF9FFFFFFFFFFFFFFFFFDFFFFFF9FFFFFFFFFF3FFFF58801CF56FCF),
    .INIT_0E(256'hFFFFFFFFFF9BFFFFFFFFFFFFFFFFFAFFFFFFCFFFFFFFFFCFFFFF6820BBFCF94F),
    .INIT_0F(256'hFFFFFFFFFF307FFFFFFFFFFFFFFFCA7FFFFFF1FFFFFFFF4FFFFFCA82435EF47B),
    .INIT_10(256'hFFFFFFFFFD067FFFFFFFFFFFFFFF887FFFFFDEFFFFFFFF3FFFFDA8098D579D99),
    .INIT_11(256'hFFFFFFFFFC207FFFFFFFFFFFFFFF0A7FFFFFFF27FFFFDAFFFFFFA0163FF75FCC),
    .INIT_12(256'hFFFFFFFFFB507FFFFFFFFFFFFFFF4A7FFFFFFF60DDD583FFFFF482DAF7FDE7D0),
    .INIT_13(256'hFFFFFFFD1694DFFFFFFFFFFFFFFFC3FFFFFFFFDE2A8A57FFFFF60141FFF5DFFE),
    .INIT_14(256'hFFFFFF708B9CDFFFFFFFFFFFFFFFFFFFFFFFFFFF7FD57FFFFFFF85A9755775FC),
    .INIT_15(256'hFFFFFFE17D3D9FFFFFFFFFFFFFFFF5557F7D7FFFFFFFFFFFFFFD5612B757F6FF),
    .INIT_16(256'hFFFFFFFFFF3D9FFFFFFFFFFFD55F5C8800A23FFFFFFFFFFFFFFFD2F6EBFFFD7F),
    .INIT_17(256'hFFFFFFFFF45E3FFFFFFFFF5778A8089777F5CB7FFFFFFFFFFFFF4BFD7EA7F73F),
    .INIT_18(256'hFFFFFFFFF2499FFFFFFFF5A822D77FFFFFFFFEBFFFFFFFFFFF67E1FFFF767DC7),
    .INIT_19(256'hFFFFFFFE3BB5CFFFFFFF003F7FFFFFFFFFFFFFCDFFFFFFFFFF07B9FFFFFF7883),
    .INIT_1A(256'hFFFFF7A37ADD67FFFFFFB7FFFFFFFFFFFFFFFF43FFFFFFFFFD3C16FFFFFFFD5F),
    .INIT_1B(256'hFFFFA2D5537FEFFFFFDF97FFFFFFFFFFFFFFFFF67FFFFFFFF431DC7FFFFFFFFF),
    .INIT_1C(256'h5595FD7FDFFDE9FFFFD71DD5A0A9DF7DFF5F7FDE9FFFFFFFF427E1BFFFFFFFFF),
    .INIT_1D(256'h55557FFFDFFF5BFFFFFDA2800AAAA0000AA08FF007FFFFFFD47FE2BFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFF71FFFFFF080A800000002A802BE227FFFFFFF8FD7B2FFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFF507FFFFF0A088A82AAA80008802009FFFFFFC8989E47FFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_016384_004 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1243,addra[14:13]}),
    .dia({open_n1247,open_n1248,open_n1249,open_n1250,open_n1251,open_n1252,open_n1253,1'b0,open_n1254}),
    .rsta(rsta),
    .doa({open_n1269,open_n1270,open_n1271,open_n1272,open_n1273,open_n1274,open_n1275,open_n1276,inst_doa_i2_004}));
  // address_offset=16384;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFEFEEE977EFFFEFF947FFF70D034C891BCFBAFFFFFFFA55561C7E1FFFFF),
    .INIT_01(256'hFFFFFFC7FFB976EFFFFFF115EFD3E407E68A2FE6BAFFFFFFF0E1561410CFFFFF),
    .INIT_02(256'hFFFFFFDBCB4D40FABFFFFF47BFE29F1CCA23FED6BBFFFFFFF0E1574D99BFFFFF),
    .INIT_03(256'hFFFFFFEF684C5B7BFFFFEF4EBFF5C7276142FFD09BFFFFFFF74156A7D8EFFFFF),
    .INIT_04(256'hFFFFFFF5FF3904CFFFFFEAFFFF949719CB9BFFC40BFFFFFFE08557A4CD6AFFFF),
    .INIT_05(256'hFFFFFFF3FDE5D423FFFFFFFFFE84D4690F53FFC013BFFFFFF0755456AA614EBF),
    .INIT_06(256'hFFFFFFFF2665554CFFFFFFFEFB5515544F1BFEE41FFFFFFFCA15556BBA1E03B5),
    .INIT_07(256'hFFFFFFFFE6185527FEFFFFFFDC555155457FFEC25FFFFFFF01555B468ADE8F84),
    .INIT_08(256'hFFFFFFFF87CB554057FFFFFF30555555556FFFF16FFFFFFF0E54591BD6EBCFFF),
    .INIT_09(256'hFFFFFFFF17A3554D6C2FFF5215555555553EFFAC7BFFFFFE945552DB875FEBFF),
    .INIT_0A(256'hFFFFFFFFF6E3555D42A8EF3355555555552BBFABFBFFFFFEB1456F8A70E7FDFF),
    .INIT_0B(256'hFFFFFFFFF0EA555553DEF1A5555555555558EFAAFFFFFFFE5155705A623FBCFB),
    .INIT_0C(256'hFFFFFFFFF8D805555053C1555555555555637BFFFFFFFFF194557A4E7B223F7F),
    .INIT_0D(256'hFFFFFFFFFD4D5555555555555555505555509EFFFFFFFFC95555D95F9DB3EF6F),
    .INIT_0E(256'hFFFFFFFFFE3E15555555555555554F5555557FFFFFFFFFAC5555888A95BA9F2F),
    .INIT_0F(256'hFFFFFFFFFE83D55555555555555562D555544EFFFFFFFF44555513FBA2FE3FB2),
    .INIT_10(256'hFFFFFFFFEF8D9555555555555555F2D55554613FFFFEFC95555359EBBBFF7E2F),
    .INIT_11(256'hFFFFFFFAB73D9555555555555555B7D5555550C7FFFFCE5555547F9FAFFB1F43),
    .INIT_12(256'hFFFFFFEF8B26C555555555555554779555555586464DFD55555B2F68AFFFBBC1),
    .INIT_13(256'hFFFFFEFAD0C63555555555555555595555555531C0386D55555B77F5FFFFA7B7),
    .INIT_14(256'hFFFFFE8E424EE555555555555555515515555505C47FD55555534E3B7FFFB0EF),
    .INIT_15(256'hFFFFFF6C8F6D25555555555555451BAE9047C55515455555555468F742FFBFBE),
    .INIT_16(256'hFFFFFFFFFDA9B555555555416FA41F1EAEFF25155555555555556AF541EAFC7B),
    .INIT_17(256'hFFFFFFBFF8DC9155555554E864D552CF0AED3ED55555555554059FFFBF3AFBAE),
    .INIT_18(256'hFFFFFFFF102B8155555416604E20FFFFFFFFF3C155555555547DB3FFFFA75DFF),
    .INIT_19(256'hFFFFFFFBA91E24555555BA18BFFFFFFFFFFFFF325555555554C91CFFFFFE5BDB),
    .INIT_1A(256'hFFFFFADBD8B2FC55555587FFFFFFFFFFFFFFFFC815555555511009FFFFFFFCAB),
    .INIT_1B(256'h5144851EC18191555565F3FFFFFFFFFFFFFFFF66D555555559A0DEFFFFFFEFFF),
    .INIT_1C(256'h54D567D01500F25555795BC8FBE97A6A55FCFF7AF5555555597FA8AFFFFFFFFF),
    .INIT_1D(256'hFFBF90013003F8555556D72AA5551FBFF45BF32ECC1555557A7FF89FFFFEBFFF),
    .INIT_1E(256'h000000000002BE555554BAAABEBAFBFFAAAEDF3AA055555558AD337FFFFFFFFF),
    .INIT_1F(256'h000000000003EE855554AAEB917D0042BAB0BAAEBB1555553590321FBFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_016384_005 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1302,addra[14:13]}),
    .dia({open_n1306,open_n1307,open_n1308,open_n1309,open_n1310,open_n1311,open_n1312,1'b0,open_n1313}),
    .rsta(rsta),
    .doa({open_n1328,open_n1329,open_n1330,open_n1331,open_n1332,open_n1333,open_n1334,open_n1335,inst_doa_i2_005}));
  // address_offset=16384;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFF045DEB8FFFFFFF2FAFFD862EF5FD1FFE2F6FFFFFFF82AAAD5DB540000),
    .INIT_01(256'hFFFFFFC554CAB6FFFFFFFEEBFFE570DF7745FFDBF3FFFFFFF8EAAA85AA140000),
    .INIT_02(256'hFFFFFFE8408ABBFFFFFFFCA3FFFD229235A8FFCFB7FFFFFFF47AAA8E43740000),
    .INIT_03(256'hFFFFFFF941CAAA7FFFFFFFFFFFEA7AC6A34BFFDE2AFFFFFFF8EAAB5D12740000),
    .INIT_04(256'hFFFFFFF0132AAABFFFFFFFFFFFBB3DBBC913FFCFBBFFFFFFE4AAAB4C06A05000),
    .INIT_05(256'hFFFFFFFE526EABFFFFFFFFFFFFEA2BB7E18FFFDFE7FFFFFFC2AAAB1923B98555),
    .INIT_06(256'hFFFFFFFE04BAAAFBFFFFFFFFFFAAAAAFA1AFFFCBE7FFFFFFFEAAAB3C62A5A6F1),
    .INIT_07(256'hFFFFFFFD81D3AABF7FFFFFFFA6AAAAAAAEAFFFFBABFFFFFFBEAAAC606B643AFB),
    .INIT_08(256'hFFFFFFFFD143AAAF0BFFFFFD1BAAAAAAAAFFFFF3DFFFFFFF1EABA92523704BFF),
    .INIT_09(256'hFFFFFFFFBCD6AAAADDAFFF81BAAAAAAAAABFFFFEFFFFFFFFBAAAAEE53A040DFF),
    .INIT_0A(256'hFFFFFFFFE612AAAABCEC040FAAAAAAAAAAC3FFFFFFFFFFFC7ABAB2002ED803BF),
    .INIT_0B(256'hFFFFFFFFEF5AAAAAABF11BFAAAAAAAAAAABFFFFFFFFFFFFEAAAAB3104DCD05BF),
    .INIT_0C(256'hFFFFFFFFF0EFAAAAAAAFFEAAAAAAAAAAAABEFFFFFFFFFFF4AAAAB9904ACF51DF),
    .INIT_0D(256'hFFFFFFFFFCBFAAAAAAAAAAAAAAAAABAAAAAFBFFFFFFFFFEFAAAAB3516311617F),
    .INIT_0E(256'hFFFFFFFFFC39EAAAAAAAAAAAAAAAA4AAAAAAB3FFFFFFFFE7AAAA94D13D42E8F3),
    .INIT_0F(256'hFFFFFFFFFEB5EAAAAAAAAAAAAAAAD5EAAAAAB9FFFFFFFF0EAAAAECC5B0077B0B),
    .INIT_10(256'hFFFFFFFFFF54AAAAAAAAAAAAAAAA40EAAAAABF7FFFFFFCFAAAAB1512F000EFDD),
    .INIT_11(256'hFFFFFFFFFA1DAAAAAAAAAAAAAAAA45EAAAAAAFAFFFFFFAEAAAAAF03A80011FF3),
    .INIT_12(256'hFFFFFFFF9CCAAAAAAAAAAAAAAAAB84EAAAAAAA8B7EF4B7AAAAAD95FA10006BEC),
    .INIT_13(256'hFFFFFFFDC71FAAAAAAAAAAAAAAAAB3AAAAAAAAB9BFA8AEAAAAAF1AAA000043F1),
    .INIT_14(256'hFFFFFFD4ADC27AAAAAAAAAAAAAAAAEAAAAAAAAABFABFAAAAAAA86ED8900013FF),
    .INIT_15(256'hFFFFFFF83F952AAAAAAAAAAAAAAAEFAEBEEFFAAAAAAAAAAAAAABFADCDC0006BE),
    .INIT_16(256'hFFFFFFFFFC80AAAAAAAAAAAABFAFA15BFEEF4BAAAAAAAAAAAAAAAEFA2844053F),
    .INIT_17(256'hFFFFFFFFFB2BFAAAAAAAABEBD0FBEA94FFFA6DAAAAAAAAAAAAFA93FEB7E1418F),
    .INIT_18(256'hFFFFFFFFCBFABEAAAAAAFD6FFF1AAFFFFFFFFAEEAAAAAAAAABBF1EFFFFD6126B),
    .INIT_19(256'hFFFFFFE78CDB5EAAAAAB7A42FFFFFFFFFFFFFF6FAAAAAAAAAA8BDCFFFFFE9ABB),
    .INIT_1A(256'hFFFFFCBDB72E2AAAAAAB9BFFFFFFFFFFFFFFFFCEEAAAAAAAAFF836BFFFFFFA02),
    .INIT_1B(256'h0550BF3A8EBE3EAAAAABCBFFFFFFFFFFFFFFFFC3AAAAAAAAA885537FFFFFFFFF),
    .INIT_1C(256'h00C15ABFEFFF36AAAAAB02F0FFEC01D01556FFD0AAAAAAAAABE115FFFFFFFFFF),
    .INIT_1D(256'hAAAABFFEFFFD4AAAAAAA8FC55555551555502F8C5AAAAAAAB3956A6FFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFC5DEAAAAA911541450400555011A15FAAAAAABE5D8DBFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFF947AAAAAA85543FFFFFBFFABE41C15AAAAAAAD1FED56FFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_016384_006 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1361,addra[14:13]}),
    .dia({open_n1365,open_n1366,open_n1367,open_n1368,open_n1369,open_n1370,open_n1371,1'b0,open_n1372}),
    .rsta(rsta),
    .doa({open_n1387,open_n1388,open_n1389,open_n1390,open_n1391,open_n1392,open_n1393,open_n1394,inst_doa_i2_006}));
  // address_offset=16384;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFCEEE3FF3FFFFFFF951FFF3CFEFFA3D2BE0FBFFFFFFFC7FFFEFD6AFFFFF),
    .INIT_01(256'hFFFFFFEEFE6BFDFFFFFFFC56FFFE9BFB8CE4FFF4FAFFFFFFFC6FFFFA17EFFFFF),
    .INIT_02(256'hFFFFFFE3EA3BFCBFFFFFFF4FFFEEB8AE9B46FFE5FEFFFFFFFCFFFFA426DFFFFF),
    .INIT_03(256'hFFFFFFF2EB7BF8FFFFFFFFEFFFFFECEADCE7FFF1A7FFFFFFF4FFFFE0B3DFFFFF),
    .INIT_04(256'hFFFFFFFFB9CBFF7FFFFFFFFFFFFEAEE6E2BBFFE147FFFFFFF7BFFFA6B79BFFFF),
    .INIT_05(256'hFFFFFFFCB8DFFF8FFFFFFFFFFFBFFFFFFBFFFFE14BFFFFFFE7FFFFA2838B6BFF),
    .INIT_06(256'hFFFFFFFDADDFFFE2FFFFFFFFFEFFFFFFFAEFFFE15BFFFFFFC2FFFE86969F495A),
    .INIT_07(256'hFFFFFFFF7DEBFFF8BFFFFFFFEFFFFFFFFFEFFFE11FFFFFFFDFFFFF8E86DFDBBF),
    .INIT_08(256'hFFFFFFFF69EFFFFFFFFFFFFAAFFFFFFFFFBFFFFC6FFFFFFFAFFFFB9B9E8BF3FF),
    .INIT_09(256'hFFFFFFFF883EFFFFF7BFFFFEFFFFFFFFFFEFFFFFFFFFFFFE3FFFFD4B9AEFE2FF),
    .INIT_0A(256'hFFFFFFFFD93EFFFFFF52EABFFFFFFFFFFFFFFFFFFFFFFFFEBFFFF87ADE6BFDBF),
    .INIT_0B(256'hFFFFFFFFE6B2FFFFFFEEAAFFFFFFFFFFFFE7FFFFFFFFFFF8FFFFF87AEE32BE7F),
    .INIT_0C(256'hFFFFFFFFFEB7FFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFABFFFF02AE861BF7F),
    .INIT_0D(256'hFFFFFFFFFFF6FFFFFFFFFFFFFFFFFEFFFFFF3FFFFFFFFFF7FFFFE5EBE9FA9FCF),
    .INIT_0E(256'hFFFFFFFFFFA3FFFFFFFFFFFFFFFFFBFFFFFFDFFFFFFFFFCFFFFFB33BF3FCF68F),
    .INIT_0F(256'hFFFFFFFFFF2EFFFFFFFFFFFFFFFFAEFFFFFFF6FFFFFFFFBFFFFFD06E9AFDF8B3),
    .INIT_10(256'hFFFFFFFFFE3FBFFFFFFFFFFFFFFFAEFFFFFFFCBFFFFFFF7FFFFF82BE0BFF6E66),
    .INIT_11(256'hFFFFFFFFFC86BFFFFFFFFFFFFFFFAAFFFFFFFF5BFFFFE0FFFFFE5AB82FFFEFC8),
    .INIT_12(256'hFFFFFFFFF7A1BFFFFFFFFFFFFFFFABFFFFFFFFA5EEEA1BFFFFFE2EA1BFFFDBE2),
    .INIT_13(256'hFFFFFFFE2969FFFFFFFFFFFFFFFFFAFFFFFFFFFF4052AFFFFFFDFF92FFFFEFFD),
    .INIT_14(256'hFFFFFFB04778FFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFEE06BFFFFAFC),
    .INIT_15(256'hFFFFFFD2BE3FAFFFFFFFFFFFFFFFFFAEBFBFFFFFFFFFFFFFFFFEF9217AFFF9FF),
    .INIT_16(256'hFFFFFFFFFF2A2FFFFFFFFFFFFFAFEEE15405EBFFFFFFFFFFFFFFE5F9D7EFFEBF),
    .INIT_17(256'hFFFFFFFFF8A17FFFFFFFFFEBBB41446FBBFAC7BFFFFFFFFFFFFFA7FEBC5BFF2F),
    .INIT_18(256'hFFFFFFFFF1866FFFFFFFFBC145EBBFFFFFFFFD2FFFFFFFFFFF9F82FFFFB9BECB),
    .INIT_19(256'hFFFFFFFC376AAFFFFFFF84FFBFFFFFFFFFFFFF9FFFFFFFFFFE7B37FFFFFFB443),
    .INIT_1A(256'hFFFFFB42A5EE8BFFFFFF2BFFFFFFFFFFFFFFFFE6FFFFFFFFFE7BA9FFFFFFFEAF),
    .INIT_1B(256'hFFFF51EAA3BFCFFFFFFF2BFFFFFFFFFFFFFFFFF8BFFFFFFFFB3EE8BFFFFFFFFF),
    .INIT_1C(256'hAA6AFEBFEFFECAFFFFFFEEEA0016EFFEEAEFBFED2FFFFFFFF95B927FFFFFFFFF),
    .INIT_1D(256'hAAAABFFFFFFFA2FFFFFE14455555551555504FF47BFFFFFFFDBFD17FFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFB7FFFFFE110000000000000017D00BFFFFFFF0F6B71FFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFEB1BFFFFE4000055555555015001012FFFFFFEB646D8BFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_016384_007 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1420,addra[14:13]}),
    .dia({open_n1424,open_n1425,open_n1426,open_n1427,open_n1428,open_n1429,open_n1430,1'b0,open_n1431}),
    .rsta(rsta),
    .doa({open_n1446,open_n1447,open_n1448,open_n1449,open_n1450,open_n1451,open_n1452,open_n1453,inst_doa_i2_007}));
  // address_offset=24576;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h555555555557F70ABEFE2FEB4000501055407EEFEBEFFFAFDE2A8AEBFFFFFFFF),
    .INIT_01(256'h55555555555FA32EBEFEBFA815555555555547BFF77FFFAEEBE6A6B3BFFFFFFF),
    .INIT_02(256'h55555555554AAA26BEFFFFA5555555555555543FA87FFFAC6AA1DD8EFFFFFFFF),
    .INIT_03(256'h55555555555FDED0AFEEBEC1555555555555551AEFBFFFA42AF1559423FFFFFF),
    .INIT_04(256'h55555555557F6EB3EFEDFE7A85555555555554D2ED4FFEA6FAF41555392FFFFF),
    .INIT_05(256'h55555555556AAAB17BEDFBABD955555555572F33A98FFF87AA9615555CD2FFFF),
    .INIT_06(256'h5555555555792AAF8AA9F9EFF1555555555DFF84FE0AFD56AAA9055555D9EFFF),
    .INIT_07(256'h5555555555BB7EAB16AA7CFBFB9555555557FFF1F94EF1CEAAA44555554CB6CB),
    .INIT_08(256'h5555555555FDFAAAC5B2EFFFFE565555756BFFF2B12AD70EAAB155555555B617),
    .INIT_09(256'h5555555555FDAAAEC32469FFFFB850004FBFFFF7BAFE189EAAF8D555555556E1),
    .INIT_0A(256'h5555555555A9BEAE57CEE4BFFFFAFFFFABFFFFAAAECD56DBABE9D55555555557),
    .INIT_0B(256'h5555555555A1EAAF1BAE7CFFFFFFFFFFFFFFFF9EECB11B9EAAA5955555555555),
    .INIT_0C(256'h5555555554BBEAAF4A7FE93FFFFFFFFFFFFFFEAEEDC73F9EAAAF055555555555),
    .INIT_0D(256'h5555555554A1AAABCFF0F55EBFFFFFFFFFFFAB0BFB3CFF9FAAB8E55555555555),
    .INIT_0E(256'h5555555550B6AAAB8FF303F4BABFFFFAAEBFECEAE073FFDBAAB7255555555555),
    .INIT_0F(256'h555555555197EAAFCFF5605201AAAAABF415EA0BEECBFFCFAAA8755555555555),
    .INIT_10(256'h5555555555FFAAAF4FFBB8FC3ABDFFABEAAD7736894FFFCFAACC355555555555),
    .INIT_11(256'h555555555406AAAF0FFC017F9655541BCA0AFEFD1C5FFF83AA9AB55555555555),
    .INIT_12(256'h55555555550AAAAB5FFD396FFFEAFFFFFFFFFFFDBD3FFF83AB44B55555555555),
    .INIT_13(256'h5555555554EEAAAB1FFF2AA7FFFFFFFFFFFFFFD23D7FFF87AF50E55555555555),
    .INIT_14(256'h555555555607AAAF1FFF2BCAFFFFFFFFFFFFFEB8E4FFFF83A855D55555555555),
    .INIT_15(256'h5555555557A2EAAE1FFFBFF20FFFFFFFFFFFEA80F1BFFF87B154955555555555),
    .INIT_16(256'h555555555484BAAE1FFFD7FED1FF903B811B5232D7FFFF9BE554055555555555),
    .INIT_17(256'h5555555555A53EAAEFFFC3E414C4055AFAA6744BD2FFFF9BC556055555555555),
    .INIT_18(256'h555555555AF55EAAEFFFE7BC87C401000157396F1FFFFF8E1556555555555555),
    .INIT_19(256'h555555555C655BAEEFFFF6F85CFB2FFE4851A3AF0FFFFFC15556955555555555),
    .INIT_1A(256'h555555555A9556FEAFFFF6EB164B5001991E60BC3FFFFFCA5556D55555555555),
    .INIT_1B(256'h555555555055557EAFFFFC6B94005202B5AA5EAF7FFFFFD25554D55555555555),
    .INIT_1C(256'h010015115F00005BEFFFFC3EC6515EFB10AB4CF4FFFFFFB15554A40510400000),
    .INIT_1D(256'h041000141A544414EFFFFEAEA8A00050A80A56BDFFFFFEF55554601500001100),
    .INIT_1E(256'h4041005408414105EFFFFF3EC1AA00AAB848BFC3FFFFFCD95556A00100440111),
    .INIT_1F(256'h5511555565941559EFFFFF4EB200000000016AE3FFFFF1D85556594545114454),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_024576_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1479,addra[14:13]}),
    .dia({open_n1483,open_n1484,open_n1485,open_n1486,open_n1487,open_n1488,open_n1489,1'b0,open_n1490}),
    .rsta(rsta),
    .doa({open_n1505,open_n1506,open_n1507,open_n1508,open_n1509,open_n1510,open_n1511,open_n1512,inst_doa_i3_000}));
  // address_offset=24576;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFF87B255554C000BFFFAFEFAABF90400155555565CC7E2BFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFF441C555544007EAAAAAAAAAAAB90006955554F5F3E5A6BFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFF514295555001AAAAAAAAAAAAAAB80029555559543BBA99FFFFFFF),
    .INIT_03(256'hFFFFFFFFFFE1F5725555003BAAAAAAAAAAAAAAE000155552556BFFBEF2FFFFFF),
    .INIT_04(256'hFFFFFFFFFFD1E549555440BAAAAAAAAAAAAAAF280165554A4576FFFFA33FFFFF),
    .INIT_05(256'hFFFFFFFFFFD50556955440EBF2AAAAAAAAA8FF8D01E5550C5540FFFFFBE6FFFF),
    .INIT_06(256'hFFFFFFFFFF859557B55142EFFEAAAAAAAAA3FFAB10A555385545EFFFFFAE9BFF),
    .INIT_07(256'hFFFFFFFFFF07D155D95242FBFC2AAAAAAAABFFFE41E550C4555BAFFFFFEB2F3F),
    .INIT_08(256'hFFFFFFFFFF47D555124B46FFFFE8AAAA8AFBFFFDC7855354555DFFFFFFFFAD3F),
    .INIT_09(256'hFFFFFFFFFF461551159E42FFFFBEFFFFEBBFFFF905D54D145518BFFFFFFFFEA9),
    .INIT_0A(256'hFFFFFFFFFF5241515567CABFFFFAFFFFABFFFFB740E02015541BBFFFFFFFFFFE),
    .INIT_0B(256'hFFFFFFFFFF5355515503E7FFFFFFFFFFFFFFFFB4018080515556BFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFF5B5551154702BFFFFFFFFFFFFFFEC901D040515551EFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFF5D5555D0164EBEBFFFFFFFFFFFABE01375005155436FFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFB495555D004285AFABFFFFAAEBFFB6407840015554E2FFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFA4D15519007F499BAFFFFFEAABE01A01DE0001555582FFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFE6D5551D0006AF9D50200015556ECB84550001555282FFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFEB55551D00122BFE6AAABFAD1BBFEFE229000595579EFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFF555559001959FFFFFFFFFFFFFFFFD4540005954AEEFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFE65555590004543FFFFFFFFFFFFFFF11600005951FBEFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFE58555190006047BFFFFFFFFFFFFF3B5500005D57FFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFED915519000040EEFFFFFFFFFFFF6D95C40005D4BFEBFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFEBF45519000011AB64015506AB57E2C500000491FFE3FFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFEAFC15540001916497AAAAFFAA9E0316500004D3FFE7FFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFF8EFE1554000044783650000002F68A54000005DBFFE6FFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFF86FF051400003458D826FFE1AA4A25590000012FFFE2FFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFA3FFC0140000555C61C8554F60A67D540000012FFFE2FFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFEFFFF8140000155E005BBEC60AA4D554000001AFFFE2FFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFF6BFFFE4000001D122500FAE40AB50510000004FFFFE0FFFEFBFFFFF),
    .INIT_1D(256'hFBEFFFFFF4EBBBFE000000112CA00000A80A28550000015FFFFE4FEEFFFFEEFF),
    .INIT_1E(256'hFFFFFFFFECFFFFFF0000007558AA00AAB80881440000026BFFFE8FFEFFBBFFFF),
    .INIT_1F(256'hFFBBFFFFEEBEBFFB100000655E0000000000E15000000A3EFFFEEBEFEFBBEEFE),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_024576_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1538,addra[14:13]}),
    .dia({open_n1542,open_n1543,open_n1544,open_n1545,open_n1546,open_n1547,open_n1548,1'b0,open_n1549}),
    .rsta(rsta),
    .doa({open_n1564,open_n1565,open_n1566,open_n1567,open_n1568,open_n1569,open_n1570,open_n1571,inst_doa_i3_001}));
  // address_offset=24576;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hAAAAAAAAAAABD1BAAAAB5555000000000000151556AAAAAA8B27C5D7FFFFFFFF),
    .INIT_01(256'hAAAAAAAAAAAFCB3AAAAB5554000000000000015551EAAAAB1F59F979FFFFFFFF),
    .INIT_02(256'hAAAAAAAAAAAFDE9EAAAA5550000000000000001554EAAAAB3FC8EE2F7FFFFFFF),
    .INIT_03(256'hAAAAAAAAAAAF4FCBAAAA5544000000000000000555EAAAA8BFD0AAEB9BFFFFFF),
    .INIT_04(256'hAAAAAAAAAABF0FF2AAAA1510400000000000000154FAAAA1FFD0AAAAFCFFFFFF),
    .INIT_05(256'hAAAAAAAAAABF3FF8EAAA15414000000000001541543AAAB7FFE1AAAAAE4BFFFF),
    .INIT_06(256'hAAAAAAAAAABE3FFD7AAF14455000000000005510453AABD2FFF4BAAAAAE47FFF),
    .INIT_07(256'hAAAAAAAAAABD3FFF3EAD15515400000000055550547AAB06FFF0BAAAAABED1EF),
    .INIT_08(256'hAAAAAAAAAAFC7FFFCBAC15555500000000115551783ABC06FFF2AAAAAAAAFB81),
    .INIT_09(256'hAAAAAAAAAAFCFFFFC2E811555515000015155551FF2AF046FFF6EAAAAAAAABFA),
    .INIT_0A(256'hAAAAAAAAAAFCFFFF80B811155550555501555515FF3BC147FFF0EAAAAAAAAAAB),
    .INIT_0B(256'hAAAAAAAAAAF8FFFF847CD4555555555555555507FE6F0547FFF8EAAAAAAAAAAA),
    .INIT_0C(256'hAAAAAAAAAAF5FFFF8518F0555555555555555447FF3D1547FFFDBAAAAAAAAAAA),
    .INIT_0D(256'hAAAAAAAAAAF2FFFF4540F004155555555555010FECC05547FFF8FAAAAAAAAAAA),
    .INIT_0E(256'hAAAAAAAAAEF3FFFF4551A551501555500415545FF8115547FFF9FAAAAAAAAAAA),
    .INIT_0F(256'hAAAAAAAAAEE3FFFF45501AA1055555555540012FF1455547FFFEBAAAAAAAAAAA),
    .INIT_10(256'hAAAAAAAAAAD7FFFF0555D6FE15000001555411BBE6855547FFEFBAAAAAAAAAAA),
    .INIT_11(256'hAAAAAAAAAB8BFFFF0554A8BFE90000056FAFFFFE8E055543FFEF7AAAAAAAAAAA),
    .INIT_12(256'hAAAAAAAAAA8FFFFF05543E3FFFFFFFFFFFFFFFFE7E155543FFBA7AAAAAAAAAAA),
    .INIT_13(256'hAAAAAAAAABDFFFFF05553FCBFFFFFFFFFFFFFFE9BC155543FFAE7AAAAAAAAAAA),
    .INIT_14(256'hAAAAAAAAABABFFFF05551BE5FFFFFFFFFFFFFFC4F8555543FEAA6AAAAAAAAAAA),
    .INIT_15(256'hAAAAAAAAAB7FFFFF05555FF12FFFFFFFFFFFFD32F0555543FAAB2AAAAAAAAAAA),
    .INIT_16(256'hAAAAAAAAAB6AFFFF05554BF55AFFEAAFEABEC1C2E1555547FAABAAAAAAAAAAAA),
    .INIT_17(256'hAAAAAAAAAA7ABFFF555543F8F040000005505FDFC1555547EAABAAAAAAAAAAAA),
    .INIT_18(256'hAAAAAAAAAF7AAFFF555553FC7C0FFFFFFFC4D71F85555547AAABAAAAAAAAAAAA),
    .INIT_19(256'hAAAAAAAAAEBAABFF555551FE3355D001F44F5D7F0555554AAAABEAAAAAAAAAAA),
    .INIT_1A(256'hAAAAAAAAADAAAAFF555551FF39F13FFF14F59D7E1555554FAAABEAAAAAAAAAAA),
    .INIT_1B(256'hAAAAAAAAA9AAAABF555554BF4FFF10054F55B1FD1555554BAAABEAAAAAAAAAAA),
    .INIT_1C(256'hAAAAAAAAADEAAAAF5555543FCDAFF001FF54B6F85555555AAAABEAAAAAAAAAAA),
    .INIT_1D(256'hAAAAAAAAAFAAAAAA5555557F935FFFFF57F5C2F45555555AAAABAAAAAAAAAAAA),
    .INIT_1E(256'hAAAAAAAAB7AAAAAA5555551FE355FF5547F75FE15555544EAAAB2AAAAAAAAAAA),
    .INIT_1F(256'hAAEEAAAAB2EBEAAE5555550FF1FFFFFFFFFF4BD55555504FAAAB2EBABAEEBBAB),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_024576_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1597,addra[14:13]}),
    .dia({open_n1601,open_n1602,open_n1603,open_n1604,open_n1605,open_n1606,open_n1607,1'b0,open_n1608}),
    .rsta(rsta),
    .doa({open_n1623,open_n1624,open_n1625,open_n1626,open_n1627,open_n1628,open_n1629,open_n1630,inst_doa_i3_002}));
  // address_offset=24576;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFF6158AAA8A02205FFFFFFFFFFDEA22AAAAAAAA90D43DBFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFA38EAAAAAA2A9FFD55FFFFFD7F402A12AAAA8D87150537FFFFFFF),
    .INIT_02(256'hFFFFFFFFFFD8299AAAAA2AA7DFFFFFFFFFFF57C8A3AAAA81C813FD9CEFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFF8FA9888A82A97FFFFFFFFFFFFFFF2AAAAAA8B08B7FF7D53FFFFFF),
    .INIT_04(256'hFFFFFFFFFFEAE0260AA2AAF0FFFFFFFFFFFFF5FCAA4AAA07A8B97FFFD39FFFFF),
    .INIT_05(256'hFFFFFFFFFF40C0ABAAA22AC35FFFFFFFFFFFDFF6284AA8322A287FFFF5F9FFFF),
    .INIT_06(256'hFFFFFFFFFFE24029C2A12147F7FFFFFFFFFDFF1D284AA96780025FFFFFD7CFFF),
    .INIT_07(256'hFFFFFFFFFF63EA0A72A32B7BD7FFFFFFFFFD7F7DA28AA1C9000DDFFFFFFD3D97),
    .INIT_08(256'hFFFFFFFFFFABE00082A3237FF5FFFFFFFDD3FF7C61EA15AB0226FFFFFFFF7C3F),
    .INIT_09(256'hFFFFFFFFFF21000000298F7FFD377555DF1FFD7E02CAFEA182A4FFFFFFFFFDD4),
    .INIT_0A(256'hFFFFFFFFFF012A002209453FFFD05FFF037FFD1182C35882828BFFFFFFFFFFFD),
    .INIT_0B(256'hFFFFFFFFFD03A8008AA9317FFFFFFF57F5FFFD1000CDC0A2000B7FFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFD2780028AA927D7FFFFFFFFF5FF5C5E0B76A0AA000A5FFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFD8E00024A810FF43FFFFFFFFFFD0B5809F0AA2880259FFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFF0C800A4AA2342FD81555500417F5BA2BC0AAA202A71FFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFF2E800ACAABFA6C755FFFF57D777CF82452AA820884BFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFF3E000ACAA235FCC2FFFFF4A0A1F47EA80AAA8A809C3FFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFF58000A4AA819FFD1FFFD77EAF5FDDD93EAAA8682347FFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFF508002EAAA6ACFFFD5FFFFFFFFFFFC00AAAA062AFD7FFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFD9200026AAA00B3FFFFFFFFFFFFF7D2ABAAAA0E8AFDDFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFD0E000A6AAA168B7FFFFFFFFFFDFD3D0A2AAA86A1FFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFF4480086AAA2AA77FFFFFFFFFFFD95E2EAAAAAE27FDBFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFD5D28086AAAAAA56902A200B54A7F7F28AAAAA68FFF1FFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFF5F6A008AAA86817CB57D5FD75C9560B0AAAAA69FFD3FFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFF4FFF8008AAAAA217D9F5FDFD7F355F82AAAAA8C7FFDBFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFC9FF6888AAAA980F7E9555D55B555224AAAAA83FFFD3FFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFF57FFDA80AAAA8887554755761F554E82AAAAA81FFFDBFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFF7FFFFE80AAAA8A8D5574D52B7D5748AAAAAAAA5FFFDBFFFFFFFFFFF),
    .INIT_1C(256'h55555F55FB5555F28AAAA868B55557F7555D5888AAAAAAA7FFFD1D5F75D55555),
    .INIT_1D(256'h5D75557D78FDDD7D8AAAAA00F55555F555557F8AAAAAAAAFFFFD157F75557F55),
    .INIT_1E(256'h555555DD76D5575F8AAAA83A2755555555D56802AAAAA9B7FFFDB55755DD7757),
    .INIT_1F(256'hFFFFFFFFD77F7FF78AAAAA980F55555555558C0AAAAAA7BFFFFDF7FFFFFFFFFD),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_024576_003 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1656,addra[14:13]}),
    .dia({open_n1660,open_n1661,open_n1662,open_n1663,open_n1664,open_n1665,open_n1666,1'b0,open_n1667}),
    .rsta(rsta),
    .doa({open_n1682,open_n1683,open_n1684,open_n1685,open_n1686,open_n1687,open_n1688,open_n1689,inst_doa_i3_003}));
  // address_offset=24576;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFF5E05FFFFF88082AAAAAAAAAAA280809FFFFFF6F39C043FFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFDEF3FFFFF0802AA800AAAAA82AAA8027FFFFF8F8EDE3C7FFFFFFF),
    .INIT_02(256'hFFFFFFFFFFF76747FFFD000A8AAAAAAAAAAA02A202FFFFD4B7C677D73FFFFFFF),
    .INIT_03(256'hFFFFFFFFFFD7ADC5DFFD80A8AAAAAAAAAAAAAA88027FFFDEF7C2FF7DE5FFFFFF),
    .INIT_04(256'hFFFFFFFFFFF7BFD95FF7000FAAAAAAAAAAAAA0AA001FFF58D7E8FFFFD6FFFFFF),
    .INIT_05(256'hFFFFFFFFFFFF9F7CFFF700BCAAAAAAAAAAAA00AA809FFD69D5D0FFFFF785FFFF),
    .INIT_06(256'hFFFFFFFFFF5F3FDC9FF40AB802AAAAAAAAAA00EA001FFC2B7FDADFFFFF5837FF),
    .INIT_07(256'hFFFFFFFFFF5EB5F727F4088422AAAAAAAAAA808A229FF4A9FFF25FFFFFF74A7F),
    .INIT_08(256'hFFFFFFFFFFDEBFFF4DF60A80082AAAAAA80C008A3CBF402BFDFBFFFFFFFF5F6A),
    .INIT_09(256'hFFFFFFFFFFDC7FFF617CA28002C2800028E00280FFBF8A2B7D717FFFFFFFFD57),
    .INIT_0A(256'hFFFFFFFFFFF4D5FFE05E2AC0002FA000FC8002C8FD9C282B7D7E7FFFFFFFFFFD),
    .INIT_0B(256'hFFFFFFFFFFF6D7FF621E6080000000A80A0002CBFD30A02BFFFC7FFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFF2FFFF60AED228000000000A00A30BFC008023FFF6DFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFF73FFFF2002708BC00000000002FC07FE8800A37FD6DFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFDD37FF7A00858AA2FEAAAAFFBE800ADF42A002BFD5C5FFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFDDB7FF7200AADDA8A0000002A828297F800002BF7755FFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFDCBFFF7A000C1F52A000000AA082275DBE0002B7F555FFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFF6FFFF7A002567FF6AAA80A3777FDFF67A000237DF79FFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFEF7FFF20023F3FFFFFFFFFFFFFFFFD3F0000A3D57D9FFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFDCDFFFF20009F6FFFFFFFFFFFFFFFDE7C0000A377FF9FFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFDF5FFF7200085DAFFFFFFFFFFFFFFE8FC00002B5FFFBFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFDB77FF720000D521FFFFFFFFFFFFC0BF000000BD7FDFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFD3FD7F720000778AD7D575FDFDD0A23F00000037FFF7FFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFD1FD5FF80002374200002AA8002A007CA00000B7FFDDFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFF59FD7FF800009DC808000000080000FC000002B7FFDDFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFF5DFF577800002FF008A00000AA0021F20000025FFFD5FFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFF47FFD5780000AF72008A0022A8002BF80000025FFFD5FFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFEFFFF57800002F7A0028288A08000FE80000025FFFD5FFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFC7FFFDD000002B7600008A2000009F60000000FFFFD5FFFDF7FFFFF),
    .INIT_1D(256'hF7DFFFFFF5D777FD0000003FC00000000000037A000000AFFFFDDFDDDFFFD5FF),
    .INIT_1E(256'hFFFFFFFFFBFFFFFF000002ADF00000000080A7D800000087FFFDFFFDFF77DFFF),
    .INIT_1F(256'hFFFFFFFFD97F7FF72000008FFA00000000009FE800000027FFFD97FFFFFFFFFD),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_024576_004 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1715,addra[14:13]}),
    .dia({open_n1719,open_n1720,open_n1721,open_n1722,open_n1723,open_n1724,open_n1725,1'b0,open_n1726}),
    .rsta(rsta),
    .doa({open_n1741,open_n1742,open_n1743,open_n1744,open_n1745,open_n1746,open_n1747,open_n1748,inst_doa_i3_004}));
  // address_offset=24576;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000000000016E0A155542AE9AAFFFAFFFFEE9ABAAC1555557F3EDEEAEFFFFFFF),
    .INIT_01(256'h00000000000EFB8515543AA2AA800AAAAA82E9EABD955544DAB7E7E6BAFFFFFF),
    .INIT_02(256'h00000000000FAE5D55553ACE8BEEBFFFAAFE022AA915552B6AD4CDDBBFBFFFFF),
    .INIT_03(256'h00000000001BCBEE2551AAB4AFAAABFEAAAEAABAFB05556C3FB4418327FFFFFF),
    .INIT_04(256'h00000000002E7FE0A55BABBA2BAAAAAAAAABA4F2BFA5558EBFB54001797FFFFF),
    .INIT_05(256'h00000000006EEBF6115AAD6EDEAAAAAAAAAB6E38ABE55602BFC710004C86FFFF),
    .INIT_06(256'h0000000001682FF9E15FABBEA6FEAAAAAEACAADA7EF45197FFA93000019DEFFF),
    .INIT_07(256'h00000000006E2FFEDC5CECBAABEFAAAAAAA6AABF3C2547DDFFB470000019F29F),
    .INIT_08(256'h0000000000FDFFFEAB1AB4EAAB2BAAAAB97EABF973548CCFFFE400000000B217),
    .INIT_09(256'h0000000000FDBFFEC8923DEAAAFC055453EAABFDEE95BDDEFFF99000000012E5),
    .INIT_0A(256'h0000000001A9ABFE0F27E9EAAAAAABFFBAAAABA1BFA7F3CBFFEC900000000007),
    .INIT_0B(256'h0000000001F0BFFF58823CEEAAAEAAAAAAAAAB96EA5F0FCFFFE4800000000000),
    .INIT_0C(256'h0000000000EABFFF0F6BEE3AAAAAAAAAAAAAAEBEAD287F8BFFFA700000000000),
    .INIT_0D(256'h0000000005F5BFFF4EBD2EDFAAAAAAAAAAAABF2EBA1EFFCEFFF5E00000000000),
    .INIT_0E(256'h0000000005F2FFFECEB70D0DBAFAAAAFFBAFB92EABB3AADAFFE6E00000000000),
    .INIT_0F(256'h000000000492FFFE8EA4613595FEAAAA8417E90AFC5AAADFFFE8300000000000),
    .INIT_10(256'h0000000004FAFFFE0EAEE9FFD5FEFFFF5502AE329C0FAADEFF8F300000000000),
    .INIT_11(256'h000000000102FFFE5FAC053FDA5003AB4F4BFAEC5E8EAAC2FF9AE00000000000),
    .INIT_12(256'h00000000015BFFFA0FAD2C7EFFBFEABFFFFFFFFF692AAAD7FE15B00000000000),
    .INIT_13(256'h0000000003AFFFFA5FAE7EF7FFFFFFFFFFFFFFF2687AAAC3FF04A00000000000),
    .INIT_14(256'h000000000312FFFE1FAB37DEBAFFFBFFFFEFFFAEE1EAAAD7FC10800000000000),
    .INIT_15(256'h0000000003AEBFFF1AABAFFB9FFFFFFFFFFFFC75E4EAAAD7E013D00000000000),
    .INIT_16(256'h000000000390AFFF1AAA96EC406EF9AAD50B3DABC3AEAADAB405400000000000),
    .INIT_17(256'h0000000000B16FFBEEAAD6EE8A7ABABF950A0E8A86EAAACE9402540000000000),
    .INIT_18(256'h000000000BB05FFBFEAAF2BB69EBFBEAAB38BEFB1AAAAADF1002000000000000),
    .INIT_19(256'h000000000C6006FEBAAAB7B9EE58FFFFE63FF96A1EAAAA900402C10100000000),
    .INIT_1A(256'h000000000A5001BEFAAAB7BE8BA8CAA8063FB9FD2AAAAA8F0402810100000000),
    .INIT_1B(256'h000000000100013EBAAAA83BBAA9AEF06F7FA1FB3AAAAA820403840010440000),
    .INIT_1C(256'h110155154BC4554FFAAAA97EDBAAE1B5EAFFBCF0EAAAABF50003940501000000),
    .INIT_1D(256'h401551045E004411BAAAABAAF6FAAAFAFEAFB3F9EAAAABE00003540511455540),
    .INIT_1E(256'h4055501459454105FAAAAB7B9BFFAAFFFE2E3BC3BAAAACD80002F51010405151),
    .INIT_1F(256'h555455542481D418EFAFFE0FB4AAAAAAAAAA0EF7FEBFF1DD5556081110441547),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_024576_005 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1774,addra[14:13]}),
    .dia({open_n1778,open_n1779,open_n1780,open_n1781,open_n1782,open_n1783,open_n1784,1'b0,open_n1785}),
    .rsta(rsta),
    .doa({open_n1800,open_n1801,open_n1802,open_n1803,open_n1804,open_n1805,open_n1806,open_n1807,inst_doa_i3_005}));
  // address_offset=24576;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFF93D2AAAAB8553BFAAAFAAAAABF40556EAAAAAF09C3E7FFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFF118FAAAABC54BEA800AAAAA82BE1555AAAAAB85F7A0A3BFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFE5151AAAAB852A8AAAAAAAAAAA039553AAAAACC073BAECDFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFE4F532AAAE5560AAAAAAAAAAAAAAE555BAAAB7056BFFBFA3FFFFFF),
    .INIT_04(256'hFFFFFFFFFFD5B15EEAAD14D12AAAAAAAAAAAA5E9556AAAEE5562BFFEE36FFFFF),
    .INIT_05(256'hFFFFFFFFFF844143AAAD13440EAAAAAAAAAB507F15AAAB8D1510BFFFBAF6FFFF),
    .INIT_06(256'hFFFFFFFFFFD18555FAAC121402AAAAAAAAAC000BC4AAAF7D5501BFFFFFEBCFFF),
    .INIT_07(256'hFFFFFFFFFFD3D5558AAC511007EAAAAAAAA4001AC1EABCD7551EFFFFFFFE3E6B),
    .INIT_08(256'hFFFFFFFFFF12C55456AA0800002BAAAAB840015F03FAF155555DFFFFFFFFAC2B),
    .INIT_09(256'hFFFFFFFFFF12155407AB4D00001110014100015B41EA08115548EFFFFFFFEEA8),
    .INIT_0A(256'hFFFFFFFFFE02155454AA8800000001550000011854ED3050554FEFFFFFFFFFFE),
    .INIT_0B(256'hFFFFFFFFFE435554406EB904000400000000010D5130C1545543BFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFE5B555445460E40000000000000047D505315145555BFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFF4D15544547CA84000000000000016053115555555F6FFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFF4C555585512EA950000000000541F147D15541555B6FFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFF1D5555C557F4DB910155500546FFF44B61554155486FFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFF3D5555C5512EFCEEFEFFFAFFEFF9B94145554555692FFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFA45555855423FFB7EFFFBB40AAFEFE301555495528FFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFF15551D55591DFFFEABFFFFFFFFFFDC415555955FEAFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFF61555195550057FFFFFFFFFFFFFFF51755554D54FEEFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFE1D555595552D03BFFFFFFFFFFFFE7F0515555D56EFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFE8C55549555115FEFFFFFFFFFFFE05D1D5555595BEFEFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFBE15549555555C77C514446FE43D7C145555594BFB2FFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFAFD550455549464DFAAFFAD00CD0607055555D7FFE7FFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFF8EFE1504555451705310000012C55A41555555CBFFE7FFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFF86FFD54455556519565555517B0519185555553FBFE3EFEFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFAFFFF5405555454811A85547F05168115555542FBFE7EFEFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFBFFFFD405555440B404FAEAE05506155555555AFBFF7FFFEFBBFFFF),
    .INIT_1C(256'hAAAAAAAAB6EEAAB145555494350000A5005504045555544FFFFF3AAABBEAAAAA),
    .INIT_1D(256'hEEBFEBBAE4FEEEAE455554002450000054056D455555555FFFFF3ABBBBEFFFEA),
    .INIT_1E(256'hAAAAAAEAF9EEAAAF4555557508550055540454015555562BFFFEDFBBBAEEBAEA),
    .INIT_1F(256'hFFFFFFFFEBBFFFFB45555565090000000001D40555555A6FFFFEFBFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_024576_006 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1833,addra[14:13]}),
    .dia({open_n1837,open_n1838,open_n1839,open_n1840,open_n1841,open_n1842,open_n1843,1'b0,open_n1844}),
    .rsta(rsta),
    .doa({open_n1859,open_n1860,open_n1861,open_n1862,open_n1863,open_n1864,open_n1865,open_n1866,inst_doa_i3_006}));
  // address_offset=24576;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFAD3EFFFFF0000000000000000100003FFFFFF9B72C083FFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFED37FFFFF4004002AA0000028010007BFFFFF3F48ED3CBFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFA9BABFFFE4010200000000000A80000BFFFFE3F99BB6B3FFFFFFF),
    .INIT_03(256'hFFFFFFFFFFEB5EDEFFFE000F000000000000000000FFFFFCFAC1FFBFDAFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFB5EA3FFFF002F8000000000000A4001AFFFE4EAD4FFFFE9FFFFFF),
    .INIT_05(256'hFFFFFFFFFFFB6EBDBFFF00BBF40000000001AFD1012FFFA2EAE0FFFFFB4AFFFF),
    .INIT_06(256'hFFFFFFFFFFAF3AAF2FFE00EBF80000000007FFF0006FFF83AAE5FFFFFFA43BFF),
    .INIT_07(256'hFFFFFFFFFFED7AAB6BFF43EFF9400000000FFFE0512FFE07AAE1BFFFFFFB85BF),
    .INIT_08(256'hFFFFFFFFFFED7AAB9EF806FFFEC1000012AFFEA0FD3FFA57AAB3FFFFFFFFAF95),
    .INIT_09(256'hFFFFFFFFFFECAAAB96B947FFFFEBEAAABAFFFEA1BF3FE117AAB2BFFFFFFFFEAB),
    .INIT_0A(256'hFFFFFFFFFFF8EAABD4EC03FFFFFFFEAAFFFFFEE7EA2A9417AAB5BFFFFFFFFFFE),
    .INIT_0B(256'hFFFFFFFFFFB9EAAB943C86FBFFFBFFFFFFFFFEF6AFEA1013AABCBFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFB1EAAB9058E4FFFFFFFFFFFFFFFB93AEA94053AAA9FFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFEB3EAABD004F43BFFFFFFFFFFFFFE8BACA10013AAACEFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFEA3AAAB5004A453AFFFFFFFFFFAAA4EBD440017AAACEFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFEE7AAAB10055EB02FAAAAAAAFF8542BB1C00017AABAAFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFEC7AAAB5000D2FB11545555001444BEE7D00017AAABAFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFF9FAAAB5001A8BFEC000050FBBBFEFF8A100013AAFB2FFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFF8EAAAF10013F2FFFFFFFFFFFFFFFFF7F400003AABE6FFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFCEAAAF10006F9BFFFFFFFFFFFFFFF9BC000013ABFF6FFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFEEAAAAB10004EE5FFFFFFFFFFFFFF81FC000003ABFF7FFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFE7FAAAB10000EA46FFFFFFFFFFFFFA2F0000007ABFF7FFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFF2FEAAB10000BB3CEFABFEBEAAE9787F0000003BFFFBFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFE2FAAAF400013BDA55555502FF43A8BC5000003AFFEAFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFA6FEAAF400006EDEA0EAAAAAA93BE4FC0000007BFFEEFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFAEFFEAB400001EE6ED3BFFFAD1AFB6F1000000AFFFEAFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFF8FFFFAB400005EB6BA16AAA85AFB87E4000001AFFFEAFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFDFFFFAB400001FF5AAA44514AFFA9ED4000001AFFFFAFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFCFBFFEE0000017B8BAAAE0BAAFFA2F90000000BFFFFBFFFEEBFFFFF),
    .INIT_1D(256'hBBEABEFFBAEBBBFE0000003FCAFAAAAAFEAF93B50000005FFFFFFFEEEEBAAABF),
    .INIT_1E(256'hFFFFFFFFB7FBFFFF0000001EF6FFAAFFFEAECBE40000004BFFFE7AEEEFBBEFBF),
    .INIT_1F(256'hFFFFFFFFE6BFFFFB1000004EF7AAAAAAAAAA3FD40000001BFFFE6BFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_024576_007 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1892,addra[14:13]}),
    .dia({open_n1896,open_n1897,open_n1898,open_n1899,open_n1900,open_n1901,open_n1902,1'b0,open_n1903}),
    .rsta(rsta),
    .doa({open_n1918,open_n1919,open_n1920,open_n1921,open_n1922,open_n1923,open_n1924,open_n1925,inst_doa_i3_007}));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i1_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_1  (
    .i0(inst_doa_i2_000),
    .i1(inst_doa_i3_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b0/B0_0 ),
    .i1(\inst_doa_mux_b0/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[0]));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_0  (
    .i0(inst_doa_i0_001),
    .i1(inst_doa_i1_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_1  (
    .i0(inst_doa_i2_001),
    .i1(inst_doa_i3_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b1/B0_0 ),
    .i1(\inst_doa_mux_b1/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[1]));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_0  (
    .i0(inst_doa_i0_002),
    .i1(inst_doa_i1_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_1  (
    .i0(inst_doa_i2_002),
    .i1(inst_doa_i3_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b2/B0_0 ),
    .i1(\inst_doa_mux_b2/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[2]));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_0  (
    .i0(inst_doa_i0_003),
    .i1(inst_doa_i1_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_1  (
    .i0(inst_doa_i2_003),
    .i1(inst_doa_i3_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b3/B0_0 ),
    .i1(\inst_doa_mux_b3/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[3]));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_0  (
    .i0(inst_doa_i0_004),
    .i1(inst_doa_i1_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_1  (
    .i0(inst_doa_i2_004),
    .i1(inst_doa_i3_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b4/B0_0 ),
    .i1(\inst_doa_mux_b4/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[4]));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_0  (
    .i0(inst_doa_i0_005),
    .i1(inst_doa_i1_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_1  (
    .i0(inst_doa_i2_005),
    .i1(inst_doa_i3_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b5/B0_0 ),
    .i1(\inst_doa_mux_b5/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[5]));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_0  (
    .i0(inst_doa_i0_006),
    .i1(inst_doa_i1_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_1  (
    .i0(inst_doa_i2_006),
    .i1(inst_doa_i3_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b6/B0_0 ),
    .i1(\inst_doa_mux_b6/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[6]));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_0  (
    .i0(inst_doa_i0_007),
    .i1(inst_doa_i1_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_1  (
    .i0(inst_doa_i2_007),
    .i1(inst_doa_i3_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b7/B0_0 ),
    .i1(\inst_doa_mux_b7/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[7]));

endmodule 

module reg_sr_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire resetout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(enout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(set),
    .q(q));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

