library verilog;
use verilog.vl_types.all;
entity ModelSim is
end ModelSim;
