library verilog;
use verilog.vl_types.all;
entity CNC_COUNTER_TB is
end CNC_COUNTER_TB;
