// Verilog netlist created by TD v4.4.433
// Wed May 15 17:41:28 2019

`timescale 1ns / 1ps
module TOP  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(1)
  (
  clk,
  i8080_CS,
  i8080_D,
  i8080_WR,
  nRST,
  LCDBK,
  LCD_B,
  LCD_CLK,
  LCD_DEN,
  LCD_G,
  LCD_HYNC,
  LCD_R,
  LCD_SYNC,
  LED,
  i8080_RS
  );

  input clk;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(3)
  input i8080_CS;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(8)
  input [7:0] i8080_D;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(12)
  input i8080_WR;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(10)
  input nRST;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(4)
  output LCDBK;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(14)
  output [7:0] LCD_B;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(21)
  output LCD_CLK;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(15)
  output LCD_DEN;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(18)
  output [7:0] LCD_G;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(20)
  output LCD_HYNC;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(16)
  output [7:0] LCD_R;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(19)
  output LCD_SYNC;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(17)
  output [1:0] LED;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(6)
  inout i8080_RS;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(9)

  wire [15:0] \D1/LineCount ;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(27)
  wire [15:0] \D1/PixelCount ;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(26)
  wire [15:0] \D1/n2 ;
  wire [15:0] \D1/n4 ;
  wire [15:0] \D1/n8 ;
  wire [15:0] \D1/n9 ;
  wire [7:0] FIFO_DI;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(55)
  wire [15:0] FIFO_DO;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(54)
  wire [7:0] LCD_B_pad;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(21)
  wire [7:0] LCD_G_pad;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(20)
  wire [7:0] LCD_R_pad;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(19)
  wire [1:0] LED_pad;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(6)
  wire [31:0] \U1/Count ;  // source/CLK_MOD.v(15)
  wire [31:0] \U1/n3 ;
  wire [31:0] \U1/n5 ;
  wire [31:0] \U2/Count ;  // source/CLK_MOD.v(15)
  wire [31:0] \U2/n3 ;
  wire [31:0] \U2/n5 ;
  wire [15:0] \U4/AddrCtrl ;  // source/LCD8080Ctrl.v(90)
  wire [4:0] \U4/LCD_Ctrl_Reg ;  // source/LCD8080Ctrl.v(43)
  wire [4:0] \U4/LCD_Pix_Reg ;  // source/LCD8080Ctrl.v(44)
  wire [15:0] \U4/n18 ;
  wire [15:0] \U4/n21 ;
  wire [7:0] i8080_D_pad;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(12)
  wire CLK_100M;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(25)
  wire \D1/FrameFlag ;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(55)
  wire \D1/add0/c0 ;
  wire \D1/add0/c1 ;
  wire \D1/add0/c10 ;
  wire \D1/add0/c11 ;
  wire \D1/add0/c12 ;
  wire \D1/add0/c13 ;
  wire \D1/add0/c14 ;
  wire \D1/add0/c15 ;
  wire \D1/add0/c2 ;
  wire \D1/add0/c3 ;
  wire \D1/add0/c4 ;
  wire \D1/add0/c5 ;
  wire \D1/add0/c6 ;
  wire \D1/add0/c7 ;
  wire \D1/add0/c8 ;
  wire \D1/add0/c9 ;
  wire \D1/add1/c0 ;
  wire \D1/add1/c1 ;
  wire \D1/add1/c10 ;
  wire \D1/add1/c11 ;
  wire \D1/add1/c12 ;
  wire \D1/add1/c13 ;
  wire \D1/add1/c14 ;
  wire \D1/add1/c15 ;
  wire \D1/add1/c2 ;
  wire \D1/add1/c3 ;
  wire \D1/add1/c4 ;
  wire \D1/add1/c5 ;
  wire \D1/add1/c6 ;
  wire \D1/add1/c7 ;
  wire \D1/add1/c8 ;
  wire \D1/add1/c9 ;
  wire \D1/lt0_c0 ;
  wire \D1/lt0_c1 ;
  wire \D1/lt0_c10 ;
  wire \D1/lt0_c11 ;
  wire \D1/lt0_c12 ;
  wire \D1/lt0_c13 ;
  wire \D1/lt0_c14 ;
  wire \D1/lt0_c15 ;
  wire \D1/lt0_c16 ;
  wire \D1/lt0_c2 ;
  wire \D1/lt0_c3 ;
  wire \D1/lt0_c4 ;
  wire \D1/lt0_c5 ;
  wire \D1/lt0_c6 ;
  wire \D1/lt0_c7 ;
  wire \D1/lt0_c8 ;
  wire \D1/lt0_c9 ;
  wire \D1/lt1_c0 ;
  wire \D1/lt1_c1 ;
  wire \D1/lt1_c10 ;
  wire \D1/lt1_c11 ;
  wire \D1/lt1_c12 ;
  wire \D1/lt1_c13 ;
  wire \D1/lt1_c14 ;
  wire \D1/lt1_c15 ;
  wire \D1/lt1_c16 ;
  wire \D1/lt1_c2 ;
  wire \D1/lt1_c3 ;
  wire \D1/lt1_c4 ;
  wire \D1/lt1_c5 ;
  wire \D1/lt1_c6 ;
  wire \D1/lt1_c7 ;
  wire \D1/lt1_c8 ;
  wire \D1/lt1_c9 ;
  wire \D1/lt2_c0 ;
  wire \D1/lt2_c1 ;
  wire \D1/lt2_c10 ;
  wire \D1/lt2_c11 ;
  wire \D1/lt2_c12 ;
  wire \D1/lt2_c13 ;
  wire \D1/lt2_c14 ;
  wire \D1/lt2_c15 ;
  wire \D1/lt2_c16 ;
  wire \D1/lt2_c2 ;
  wire \D1/lt2_c3 ;
  wire \D1/lt2_c4 ;
  wire \D1/lt2_c5 ;
  wire \D1/lt2_c6 ;
  wire \D1/lt2_c7 ;
  wire \D1/lt2_c8 ;
  wire \D1/lt2_c9 ;
  wire \D1/lt3_c0 ;
  wire \D1/lt3_c1 ;
  wire \D1/lt3_c10 ;
  wire \D1/lt3_c11 ;
  wire \D1/lt3_c12 ;
  wire \D1/lt3_c13 ;
  wire \D1/lt3_c14 ;
  wire \D1/lt3_c15 ;
  wire \D1/lt3_c16 ;
  wire \D1/lt3_c2 ;
  wire \D1/lt3_c3 ;
  wire \D1/lt3_c4 ;
  wire \D1/lt3_c5 ;
  wire \D1/lt3_c6 ;
  wire \D1/lt3_c7 ;
  wire \D1/lt3_c8 ;
  wire \D1/lt3_c9 ;
  wire \D1/lt4_c0 ;
  wire \D1/lt4_c1 ;
  wire \D1/lt4_c10 ;
  wire \D1/lt4_c11 ;
  wire \D1/lt4_c12 ;
  wire \D1/lt4_c13 ;
  wire \D1/lt4_c14 ;
  wire \D1/lt4_c15 ;
  wire \D1/lt4_c16 ;
  wire \D1/lt4_c2 ;
  wire \D1/lt4_c3 ;
  wire \D1/lt4_c4 ;
  wire \D1/lt4_c5 ;
  wire \D1/lt4_c6 ;
  wire \D1/lt4_c7 ;
  wire \D1/lt4_c8 ;
  wire \D1/lt4_c9 ;
  wire \D1/lt5_c0 ;
  wire \D1/lt5_c1 ;
  wire \D1/lt5_c10 ;
  wire \D1/lt5_c11 ;
  wire \D1/lt5_c12 ;
  wire \D1/lt5_c13 ;
  wire \D1/lt5_c14 ;
  wire \D1/lt5_c15 ;
  wire \D1/lt5_c16 ;
  wire \D1/lt5_c2 ;
  wire \D1/lt5_c3 ;
  wire \D1/lt5_c4 ;
  wire \D1/lt5_c5 ;
  wire \D1/lt5_c6 ;
  wire \D1/lt5_c7 ;
  wire \D1/lt5_c8 ;
  wire \D1/lt5_c9 ;
  wire \D1/lt6_c0 ;
  wire \D1/lt6_c1 ;
  wire \D1/lt6_c10 ;
  wire \D1/lt6_c11 ;
  wire \D1/lt6_c12 ;
  wire \D1/lt6_c13 ;
  wire \D1/lt6_c14 ;
  wire \D1/lt6_c15 ;
  wire \D1/lt6_c16 ;
  wire \D1/lt6_c2 ;
  wire \D1/lt6_c3 ;
  wire \D1/lt6_c4 ;
  wire \D1/lt6_c5 ;
  wire \D1/lt6_c6 ;
  wire \D1/lt6_c7 ;
  wire \D1/lt6_c8 ;
  wire \D1/lt6_c9 ;
  wire \D1/lt7_c0 ;
  wire \D1/lt7_c1 ;
  wire \D1/lt7_c10 ;
  wire \D1/lt7_c11 ;
  wire \D1/lt7_c12 ;
  wire \D1/lt7_c13 ;
  wire \D1/lt7_c14 ;
  wire \D1/lt7_c15 ;
  wire \D1/lt7_c16 ;
  wire \D1/lt7_c2 ;
  wire \D1/lt7_c3 ;
  wire \D1/lt7_c4 ;
  wire \D1/lt7_c5 ;
  wire \D1/lt7_c6 ;
  wire \D1/lt7_c7 ;
  wire \D1/lt7_c8 ;
  wire \D1/lt7_c9 ;
  wire \D1/lt8_c0 ;
  wire \D1/lt8_c1 ;
  wire \D1/lt8_c10 ;
  wire \D1/lt8_c11 ;
  wire \D1/lt8_c12 ;
  wire \D1/lt8_c13 ;
  wire \D1/lt8_c14 ;
  wire \D1/lt8_c15 ;
  wire \D1/lt8_c16 ;
  wire \D1/lt8_c2 ;
  wire \D1/lt8_c3 ;
  wire \D1/lt8_c4 ;
  wire \D1/lt8_c5 ;
  wire \D1/lt8_c6 ;
  wire \D1/lt8_c7 ;
  wire \D1/lt8_c8 ;
  wire \D1/lt8_c9 ;
  wire \D1/lt9_c0 ;
  wire \D1/lt9_c1 ;
  wire \D1/lt9_c10 ;
  wire \D1/lt9_c11 ;
  wire \D1/lt9_c12 ;
  wire \D1/lt9_c13 ;
  wire \D1/lt9_c14 ;
  wire \D1/lt9_c15 ;
  wire \D1/lt9_c16 ;
  wire \D1/lt9_c2 ;
  wire \D1/lt9_c3 ;
  wire \D1/lt9_c4 ;
  wire \D1/lt9_c5 ;
  wire \D1/lt9_c6 ;
  wire \D1/lt9_c7 ;
  wire \D1/lt9_c8 ;
  wire \D1/lt9_c9 ;
  wire \D1/mux3_b0_sel_is_0_o ;
  wire \D1/n13 ;
  wire \D1/n14 ;
  wire \D1/n15 ;
  wire \D1/n17 ;
  wire \D1/n18 ;
  wire \D1/n20 ;
  wire \D1/n22 ;
  wire \D1/n24 ;
  wire \D1/n26 ;
  wire \D1/n28 ;
  wire \FIFO0/logic_fifo_full ;
  wire \FIFO0/logic_fifo_full_neg ;
  wire FIFO_CLK_W;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(49)
  wire FIFO_EMPTY;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(52)
  wire FIFO_RE;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(50)
  wire FIFO_RST;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(47)
  wire FIFO_WE;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(51)
  wire LCD_CLK_pad;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(15)
  wire LCD_DEN_pad;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(18)
  wire LCD_HYNC_pad;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(16)
  wire LCD_SYNC_pad;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(17)
  wire \PLL1/clk0_buf ;  // al_ip/LCDPLL.v(39)
  wire \U1/add0/c0 ;
  wire \U1/add0/c1 ;
  wire \U1/add0/c10 ;
  wire \U1/add0/c11 ;
  wire \U1/add0/c12 ;
  wire \U1/add0/c13 ;
  wire \U1/add0/c14 ;
  wire \U1/add0/c15 ;
  wire \U1/add0/c16 ;
  wire \U1/add0/c17 ;
  wire \U1/add0/c18 ;
  wire \U1/add0/c19 ;
  wire \U1/add0/c2 ;
  wire \U1/add0/c20 ;
  wire \U1/add0/c21 ;
  wire \U1/add0/c22 ;
  wire \U1/add0/c23 ;
  wire \U1/add0/c24 ;
  wire \U1/add0/c25 ;
  wire \U1/add0/c26 ;
  wire \U1/add0/c27 ;
  wire \U1/add0/c28 ;
  wire \U1/add0/c29 ;
  wire \U1/add0/c3 ;
  wire \U1/add0/c30 ;
  wire \U1/add0/c31 ;
  wire \U1/add0/c4 ;
  wire \U1/add0/c5 ;
  wire \U1/add0/c6 ;
  wire \U1/add0/c7 ;
  wire \U1/add0/c8 ;
  wire \U1/add0/c9 ;
  wire \U1/n1 ;
  wire \U1/n2 ;
  wire \U2/add0/c0 ;
  wire \U2/add0/c1 ;
  wire \U2/add0/c10 ;
  wire \U2/add0/c11 ;
  wire \U2/add0/c12 ;
  wire \U2/add0/c13 ;
  wire \U2/add0/c14 ;
  wire \U2/add0/c15 ;
  wire \U2/add0/c16 ;
  wire \U2/add0/c17 ;
  wire \U2/add0/c18 ;
  wire \U2/add0/c19 ;
  wire \U2/add0/c2 ;
  wire \U2/add0/c20 ;
  wire \U2/add0/c21 ;
  wire \U2/add0/c22 ;
  wire \U2/add0/c23 ;
  wire \U2/add0/c24 ;
  wire \U2/add0/c25 ;
  wire \U2/add0/c26 ;
  wire \U2/add0/c27 ;
  wire \U2/add0/c28 ;
  wire \U2/add0/c29 ;
  wire \U2/add0/c3 ;
  wire \U2/add0/c30 ;
  wire \U2/add0/c31 ;
  wire \U2/add0/c4 ;
  wire \U2/add0/c5 ;
  wire \U2/add0/c6 ;
  wire \U2/add0/c7 ;
  wire \U2/add0/c8 ;
  wire \U2/add0/c9 ;
  wire \U2/n1 ;
  wire \U2/n2 ;
  wire \U4/FrameSync ;  // source/LCD8080Ctrl.v(54)
  wire \U4/add0/c0 ;
  wire \U4/add0/c1 ;
  wire \U4/add0/c10 ;
  wire \U4/add0/c11 ;
  wire \U4/add0/c12 ;
  wire \U4/add0/c13 ;
  wire \U4/add0/c14 ;
  wire \U4/add0/c15 ;
  wire \U4/add0/c2 ;
  wire \U4/add0/c3 ;
  wire \U4/add0/c4 ;
  wire \U4/add0/c5 ;
  wire \U4/add0/c6 ;
  wire \U4/add0/c7 ;
  wire \U4/add0/c8 ;
  wire \U4/add0/c9 ;
  wire \U4/lt0_c0 ;
  wire \U4/lt0_c1 ;
  wire \U4/lt0_c10 ;
  wire \U4/lt0_c11 ;
  wire \U4/lt0_c12 ;
  wire \U4/lt0_c13 ;
  wire \U4/lt0_c14 ;
  wire \U4/lt0_c15 ;
  wire \U4/lt0_c16 ;
  wire \U4/lt0_c2 ;
  wire \U4/lt0_c3 ;
  wire \U4/lt0_c4 ;
  wire \U4/lt0_c5 ;
  wire \U4/lt0_c6 ;
  wire \U4/lt0_c7 ;
  wire \U4/lt0_c8 ;
  wire \U4/lt0_c9 ;
  wire \U4/lt1_c0 ;
  wire \U4/lt1_c1 ;
  wire \U4/lt1_c10 ;
  wire \U4/lt1_c11 ;
  wire \U4/lt1_c12 ;
  wire \U4/lt1_c13 ;
  wire \U4/lt1_c14 ;
  wire \U4/lt1_c15 ;
  wire \U4/lt1_c16 ;
  wire \U4/lt1_c2 ;
  wire \U4/lt1_c3 ;
  wire \U4/lt1_c4 ;
  wire \U4/lt1_c5 ;
  wire \U4/lt1_c6 ;
  wire \U4/lt1_c7 ;
  wire \U4/lt1_c8 ;
  wire \U4/lt1_c9 ;
  wire \U4/lt2_c0 ;
  wire \U4/lt2_c1 ;
  wire \U4/lt2_c10 ;
  wire \U4/lt2_c11 ;
  wire \U4/lt2_c12 ;
  wire \U4/lt2_c13 ;
  wire \U4/lt2_c14 ;
  wire \U4/lt2_c15 ;
  wire \U4/lt2_c16 ;
  wire \U4/lt2_c2 ;
  wire \U4/lt2_c3 ;
  wire \U4/lt2_c4 ;
  wire \U4/lt2_c5 ;
  wire \U4/lt2_c6 ;
  wire \U4/lt2_c7 ;
  wire \U4/lt2_c8 ;
  wire \U4/lt2_c9 ;
  wire \U4/lt3_c0 ;
  wire \U4/lt3_c1 ;
  wire \U4/lt3_c10 ;
  wire \U4/lt3_c11 ;
  wire \U4/lt3_c12 ;
  wire \U4/lt3_c13 ;
  wire \U4/lt3_c14 ;
  wire \U4/lt3_c15 ;
  wire \U4/lt3_c16 ;
  wire \U4/lt3_c2 ;
  wire \U4/lt3_c3 ;
  wire \U4/lt3_c4 ;
  wire \U4/lt3_c5 ;
  wire \U4/lt3_c6 ;
  wire \U4/lt3_c7 ;
  wire \U4/lt3_c8 ;
  wire \U4/lt3_c9 ;
  wire \U4/lt4_c0 ;
  wire \U4/lt4_c1 ;
  wire \U4/lt4_c10 ;
  wire \U4/lt4_c11 ;
  wire \U4/lt4_c12 ;
  wire \U4/lt4_c13 ;
  wire \U4/lt4_c14 ;
  wire \U4/lt4_c15 ;
  wire \U4/lt4_c16 ;
  wire \U4/lt4_c2 ;
  wire \U4/lt4_c3 ;
  wire \U4/lt4_c4 ;
  wire \U4/lt4_c5 ;
  wire \U4/lt4_c6 ;
  wire \U4/lt4_c7 ;
  wire \U4/lt4_c8 ;
  wire \U4/lt4_c9 ;
  wire \U4/lt5_c0 ;
  wire \U4/lt5_c1 ;
  wire \U4/lt5_c10 ;
  wire \U4/lt5_c11 ;
  wire \U4/lt5_c12 ;
  wire \U4/lt5_c13 ;
  wire \U4/lt5_c14 ;
  wire \U4/lt5_c15 ;
  wire \U4/lt5_c16 ;
  wire \U4/lt5_c2 ;
  wire \U4/lt5_c3 ;
  wire \U4/lt5_c4 ;
  wire \U4/lt5_c5 ;
  wire \U4/lt5_c6 ;
  wire \U4/lt5_c7 ;
  wire \U4/lt5_c8 ;
  wire \U4/lt5_c9 ;
  wire \U4/lt6_c0 ;
  wire \U4/lt6_c1 ;
  wire \U4/lt6_c10 ;
  wire \U4/lt6_c11 ;
  wire \U4/lt6_c12 ;
  wire \U4/lt6_c13 ;
  wire \U4/lt6_c14 ;
  wire \U4/lt6_c15 ;
  wire \U4/lt6_c16 ;
  wire \U4/lt6_c2 ;
  wire \U4/lt6_c3 ;
  wire \U4/lt6_c4 ;
  wire \U4/lt6_c5 ;
  wire \U4/lt6_c6 ;
  wire \U4/lt6_c7 ;
  wire \U4/lt6_c8 ;
  wire \U4/lt6_c9 ;
  wire \U4/lt7_c0 ;
  wire \U4/lt7_c1 ;
  wire \U4/lt7_c10 ;
  wire \U4/lt7_c11 ;
  wire \U4/lt7_c12 ;
  wire \U4/lt7_c13 ;
  wire \U4/lt7_c14 ;
  wire \U4/lt7_c15 ;
  wire \U4/lt7_c16 ;
  wire \U4/lt7_c2 ;
  wire \U4/lt7_c3 ;
  wire \U4/lt7_c4 ;
  wire \U4/lt7_c5 ;
  wire \U4/lt7_c6 ;
  wire \U4/lt7_c7 ;
  wire \U4/lt7_c8 ;
  wire \U4/lt7_c9 ;
  wire \U4/mux0_b3_sel_is_3_o ;
  wire \U4/mux10_b0_sel_is_0_o ;
  wire \U4/mux1_b0_sel_is_3_o ;
  wire \U4/mux2_b0_sel_is_3_o ;
  wire \U4/n17 ;
  wire \U4/n23 ;
  wire \U4/n27 ;
  wire \U4/n31 ;
  wire \U4/n33 ;
  wire \U4/n37 ;
  wire \U4/n39 ;
  wire \U4/n43 ;
  wire _al_u125_o;
  wire _al_u149_o;
  wire _al_u150_o;
  wire _al_u151_o;
  wire _al_u152_o;
  wire _al_u153_o;
  wire _al_u155_o;
  wire _al_u156_o;
  wire _al_u157_o;
  wire _al_u158_o;
  wire _al_u159_o;
  wire _al_u160_o;
  wire _al_u161_o;
  wire _al_u162_o;
  wire _al_u164_o;
  wire _al_u165_o;
  wire _al_u166_o;
  wire _al_u167_o;
  wire _al_u168_o;
  wire _al_u169_o;
  wire _al_u170_o;
  wire _al_u171_o;
  wire _al_u173_o;
  wire _al_u174_o;
  wire _al_u175_o;
  wire _al_u176_o;
  wire _al_u177_o;
  wire _al_u276_o;
  wire _al_u277_o;
  wire _al_u278_o;
  wire _al_u279_o;
  wire _al_u283_o;
  wire _al_u287_o;
  wire _al_u288_o;
  wire clk_pad;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(3)
  wire i8080_CS_pad;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(8)
  wire i8080_RS_pad;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(9)
  wire i8080_WR_pad;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(10)
  wire nRST_pad;  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(4)

  reg_ar_as_w1 \D1/FrameFlag_reg  (
    .clk(LCD_CLK_pad),
    .d(\D1/n13 ),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/FrameFlag ));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(84)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add0/u0  (
    .a(\D1/LineCount [0]),
    .b(1'b1),
    .c(\D1/add0/c0 ),
    .o({\D1/add0/c1 ,\D1/n2 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add0/u1  (
    .a(\D1/LineCount [1]),
    .b(1'b0),
    .c(\D1/add0/c1 ),
    .o({\D1/add0/c2 ,\D1/n2 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add0/u10  (
    .a(\D1/LineCount [10]),
    .b(1'b0),
    .c(\D1/add0/c10 ),
    .o({\D1/add0/c11 ,\D1/n2 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add0/u11  (
    .a(\D1/LineCount [11]),
    .b(1'b0),
    .c(\D1/add0/c11 ),
    .o({\D1/add0/c12 ,\D1/n2 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add0/u12  (
    .a(\D1/LineCount [12]),
    .b(1'b0),
    .c(\D1/add0/c12 ),
    .o({\D1/add0/c13 ,\D1/n2 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add0/u13  (
    .a(\D1/LineCount [13]),
    .b(1'b0),
    .c(\D1/add0/c13 ),
    .o({\D1/add0/c14 ,\D1/n2 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add0/u14  (
    .a(\D1/LineCount [14]),
    .b(1'b0),
    .c(\D1/add0/c14 ),
    .o({\D1/add0/c15 ,\D1/n2 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add0/u15  (
    .a(\D1/LineCount [15]),
    .b(1'b0),
    .c(\D1/add0/c15 ),
    .o({open_n0,\D1/n2 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add0/u2  (
    .a(\D1/LineCount [2]),
    .b(1'b0),
    .c(\D1/add0/c2 ),
    .o({\D1/add0/c3 ,\D1/n2 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add0/u3  (
    .a(\D1/LineCount [3]),
    .b(1'b0),
    .c(\D1/add0/c3 ),
    .o({\D1/add0/c4 ,\D1/n2 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add0/u4  (
    .a(\D1/LineCount [4]),
    .b(1'b0),
    .c(\D1/add0/c4 ),
    .o({\D1/add0/c5 ,\D1/n2 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add0/u5  (
    .a(\D1/LineCount [5]),
    .b(1'b0),
    .c(\D1/add0/c5 ),
    .o({\D1/add0/c6 ,\D1/n2 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add0/u6  (
    .a(\D1/LineCount [6]),
    .b(1'b0),
    .c(\D1/add0/c6 ),
    .o({\D1/add0/c7 ,\D1/n2 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add0/u7  (
    .a(\D1/LineCount [7]),
    .b(1'b0),
    .c(\D1/add0/c7 ),
    .o({\D1/add0/c8 ,\D1/n2 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add0/u8  (
    .a(\D1/LineCount [8]),
    .b(1'b0),
    .c(\D1/add0/c8 ),
    .o({\D1/add0/c9 ,\D1/n2 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add0/u9  (
    .a(\D1/LineCount [9]),
    .b(1'b0),
    .c(\D1/add0/c9 ),
    .o({\D1/add0/c10 ,\D1/n2 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \D1/add0/ucin  (
    .a(1'b0),
    .o({\D1/add0/c0 ,open_n3}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add1/u0  (
    .a(\D1/PixelCount [0]),
    .b(1'b1),
    .c(\D1/add1/c0 ),
    .o({\D1/add1/c1 ,\D1/n4 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add1/u1  (
    .a(\D1/PixelCount [1]),
    .b(1'b0),
    .c(\D1/add1/c1 ),
    .o({\D1/add1/c2 ,\D1/n4 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add1/u10  (
    .a(\D1/PixelCount [10]),
    .b(1'b0),
    .c(\D1/add1/c10 ),
    .o({\D1/add1/c11 ,\D1/n4 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add1/u11  (
    .a(\D1/PixelCount [11]),
    .b(1'b0),
    .c(\D1/add1/c11 ),
    .o({\D1/add1/c12 ,\D1/n4 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add1/u12  (
    .a(\D1/PixelCount [12]),
    .b(1'b0),
    .c(\D1/add1/c12 ),
    .o({\D1/add1/c13 ,\D1/n4 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add1/u13  (
    .a(\D1/PixelCount [13]),
    .b(1'b0),
    .c(\D1/add1/c13 ),
    .o({\D1/add1/c14 ,\D1/n4 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add1/u14  (
    .a(\D1/PixelCount [14]),
    .b(1'b0),
    .c(\D1/add1/c14 ),
    .o({\D1/add1/c15 ,\D1/n4 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add1/u15  (
    .a(\D1/PixelCount [15]),
    .b(1'b0),
    .c(\D1/add1/c15 ),
    .o({open_n4,\D1/n4 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add1/u2  (
    .a(\D1/PixelCount [2]),
    .b(1'b0),
    .c(\D1/add1/c2 ),
    .o({\D1/add1/c3 ,\D1/n4 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add1/u3  (
    .a(\D1/PixelCount [3]),
    .b(1'b0),
    .c(\D1/add1/c3 ),
    .o({\D1/add1/c4 ,\D1/n4 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add1/u4  (
    .a(\D1/PixelCount [4]),
    .b(1'b0),
    .c(\D1/add1/c4 ),
    .o({\D1/add1/c5 ,\D1/n4 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add1/u5  (
    .a(\D1/PixelCount [5]),
    .b(1'b0),
    .c(\D1/add1/c5 ),
    .o({\D1/add1/c6 ,\D1/n4 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add1/u6  (
    .a(\D1/PixelCount [6]),
    .b(1'b0),
    .c(\D1/add1/c6 ),
    .o({\D1/add1/c7 ,\D1/n4 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add1/u7  (
    .a(\D1/PixelCount [7]),
    .b(1'b0),
    .c(\D1/add1/c7 ),
    .o({\D1/add1/c8 ,\D1/n4 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add1/u8  (
    .a(\D1/PixelCount [8]),
    .b(1'b0),
    .c(\D1/add1/c8 ),
    .o({\D1/add1/c9 ,\D1/n4 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \D1/add1/u9  (
    .a(\D1/PixelCount [9]),
    .b(1'b0),
    .c(\D1/add1/c9 ),
    .o({\D1/add1/c10 ,\D1/n4 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \D1/add1/ucin  (
    .a(1'b0),
    .o({\D1/add1/c0 ,open_n7}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt0_0  (
    .a(1'b0),
    .b(\D1/PixelCount [0]),
    .c(\D1/lt0_c0 ),
    .o({\D1/lt0_c1 ,open_n8}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt0_1  (
    .a(1'b0),
    .b(\D1/PixelCount [1]),
    .c(\D1/lt0_c1 ),
    .o({\D1/lt0_c2 ,open_n9}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt0_10  (
    .a(1'b0),
    .b(\D1/PixelCount [10]),
    .c(\D1/lt0_c10 ),
    .o({\D1/lt0_c11 ,open_n10}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt0_11  (
    .a(1'b0),
    .b(\D1/PixelCount [11]),
    .c(\D1/lt0_c11 ),
    .o({\D1/lt0_c12 ,open_n11}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt0_12  (
    .a(1'b0),
    .b(\D1/PixelCount [12]),
    .c(\D1/lt0_c12 ),
    .o({\D1/lt0_c13 ,open_n12}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt0_13  (
    .a(1'b0),
    .b(\D1/PixelCount [13]),
    .c(\D1/lt0_c13 ),
    .o({\D1/lt0_c14 ,open_n13}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt0_14  (
    .a(1'b0),
    .b(\D1/PixelCount [14]),
    .c(\D1/lt0_c14 ),
    .o({\D1/lt0_c15 ,open_n14}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt0_15  (
    .a(1'b0),
    .b(\D1/PixelCount [15]),
    .c(\D1/lt0_c15 ),
    .o({\D1/lt0_c16 ,open_n15}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt0_2  (
    .a(1'b1),
    .b(\D1/PixelCount [2]),
    .c(\D1/lt0_c2 ),
    .o({\D1/lt0_c3 ,open_n16}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt0_3  (
    .a(1'b0),
    .b(\D1/PixelCount [3]),
    .c(\D1/lt0_c3 ),
    .o({\D1/lt0_c4 ,open_n17}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt0_4  (
    .a(1'b1),
    .b(\D1/PixelCount [4]),
    .c(\D1/lt0_c4 ),
    .o({\D1/lt0_c5 ,open_n18}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt0_5  (
    .a(1'b0),
    .b(\D1/PixelCount [5]),
    .c(\D1/lt0_c5 ),
    .o({\D1/lt0_c6 ,open_n19}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt0_6  (
    .a(1'b0),
    .b(\D1/PixelCount [6]),
    .c(\D1/lt0_c6 ),
    .o({\D1/lt0_c7 ,open_n20}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt0_7  (
    .a(1'b0),
    .b(\D1/PixelCount [7]),
    .c(\D1/lt0_c7 ),
    .o({\D1/lt0_c8 ,open_n21}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt0_8  (
    .a(1'b0),
    .b(\D1/PixelCount [8]),
    .c(\D1/lt0_c8 ),
    .o({\D1/lt0_c9 ,open_n22}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt0_9  (
    .a(1'b0),
    .b(\D1/PixelCount [9]),
    .c(\D1/lt0_c9 ),
    .o({\D1/lt0_c10 ,open_n23}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \D1/lt0_cin  (
    .a(1'b1),
    .o({\D1/lt0_c0 ,open_n26}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt0_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\D1/lt0_c16 ),
    .o({open_n27,\D1/n14 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt1_0  (
    .a(\D1/PixelCount [0]),
    .b(1'b1),
    .c(\D1/lt1_c0 ),
    .o({\D1/lt1_c1 ,open_n28}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt1_1  (
    .a(\D1/PixelCount [1]),
    .b(1'b1),
    .c(\D1/lt1_c1 ),
    .o({\D1/lt1_c2 ,open_n29}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt1_10  (
    .a(\D1/PixelCount [10]),
    .b(1'b0),
    .c(\D1/lt1_c10 ),
    .o({\D1/lt1_c11 ,open_n30}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt1_11  (
    .a(\D1/PixelCount [11]),
    .b(1'b0),
    .c(\D1/lt1_c11 ),
    .o({\D1/lt1_c12 ,open_n31}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt1_12  (
    .a(\D1/PixelCount [12]),
    .b(1'b0),
    .c(\D1/lt1_c12 ),
    .o({\D1/lt1_c13 ,open_n32}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt1_13  (
    .a(\D1/PixelCount [13]),
    .b(1'b0),
    .c(\D1/lt1_c13 ),
    .o({\D1/lt1_c14 ,open_n33}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt1_14  (
    .a(\D1/PixelCount [14]),
    .b(1'b0),
    .c(\D1/lt1_c14 ),
    .o({\D1/lt1_c15 ,open_n34}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt1_15  (
    .a(\D1/PixelCount [15]),
    .b(1'b0),
    .c(\D1/lt1_c15 ),
    .o({\D1/lt1_c16 ,open_n35}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt1_2  (
    .a(\D1/PixelCount [2]),
    .b(1'b1),
    .c(\D1/lt1_c2 ),
    .o({\D1/lt1_c3 ,open_n36}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt1_3  (
    .a(\D1/PixelCount [3]),
    .b(1'b1),
    .c(\D1/lt1_c3 ),
    .o({\D1/lt1_c4 ,open_n37}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt1_4  (
    .a(\D1/PixelCount [4]),
    .b(1'b0),
    .c(\D1/lt1_c4 ),
    .o({\D1/lt1_c5 ,open_n38}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt1_5  (
    .a(\D1/PixelCount [5]),
    .b(1'b0),
    .c(\D1/lt1_c5 ),
    .o({\D1/lt1_c6 ,open_n39}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt1_6  (
    .a(\D1/PixelCount [6]),
    .b(1'b1),
    .c(\D1/lt1_c6 ),
    .o({\D1/lt1_c7 ,open_n40}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt1_7  (
    .a(\D1/PixelCount [7]),
    .b(1'b1),
    .c(\D1/lt1_c7 ),
    .o({\D1/lt1_c8 ,open_n41}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt1_8  (
    .a(\D1/PixelCount [8]),
    .b(1'b0),
    .c(\D1/lt1_c8 ),
    .o({\D1/lt1_c9 ,open_n42}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt1_9  (
    .a(\D1/PixelCount [9]),
    .b(1'b1),
    .c(\D1/lt1_c9 ),
    .o({\D1/lt1_c10 ,open_n43}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \D1/lt1_cin  (
    .a(1'b0),
    .o({\D1/lt1_c0 ,open_n46}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt1_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\D1/lt1_c16 ),
    .o({open_n47,\D1/n15 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt2_0  (
    .a(\D1/LineCount [0]),
    .b(1'b0),
    .c(\D1/lt2_c0 ),
    .o({\D1/lt2_c1 ,open_n48}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt2_1  (
    .a(\D1/LineCount [1]),
    .b(1'b1),
    .c(\D1/lt2_c1 ),
    .o({\D1/lt2_c2 ,open_n49}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt2_10  (
    .a(\D1/LineCount [10]),
    .b(1'b0),
    .c(\D1/lt2_c10 ),
    .o({\D1/lt2_c11 ,open_n50}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt2_11  (
    .a(\D1/LineCount [11]),
    .b(1'b0),
    .c(\D1/lt2_c11 ),
    .o({\D1/lt2_c12 ,open_n51}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt2_12  (
    .a(\D1/LineCount [12]),
    .b(1'b0),
    .c(\D1/lt2_c12 ),
    .o({\D1/lt2_c13 ,open_n52}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt2_13  (
    .a(\D1/LineCount [13]),
    .b(1'b0),
    .c(\D1/lt2_c13 ),
    .o({\D1/lt2_c14 ,open_n53}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt2_14  (
    .a(\D1/LineCount [14]),
    .b(1'b0),
    .c(\D1/lt2_c14 ),
    .o({\D1/lt2_c15 ,open_n54}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt2_15  (
    .a(\D1/LineCount [15]),
    .b(1'b0),
    .c(\D1/lt2_c15 ),
    .o({\D1/lt2_c16 ,open_n55}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt2_2  (
    .a(\D1/LineCount [2]),
    .b(1'b0),
    .c(\D1/lt2_c2 ),
    .o({\D1/lt2_c3 ,open_n56}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt2_3  (
    .a(\D1/LineCount [3]),
    .b(1'b1),
    .c(\D1/lt2_c3 ),
    .o({\D1/lt2_c4 ,open_n57}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt2_4  (
    .a(\D1/LineCount [4]),
    .b(1'b0),
    .c(\D1/lt2_c4 ),
    .o({\D1/lt2_c5 ,open_n58}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt2_5  (
    .a(\D1/LineCount [5]),
    .b(1'b0),
    .c(\D1/lt2_c5 ),
    .o({\D1/lt2_c6 ,open_n59}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt2_6  (
    .a(\D1/LineCount [6]),
    .b(1'b0),
    .c(\D1/lt2_c6 ),
    .o({\D1/lt2_c7 ,open_n60}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt2_7  (
    .a(\D1/LineCount [7]),
    .b(1'b0),
    .c(\D1/lt2_c7 ),
    .o({\D1/lt2_c8 ,open_n61}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt2_8  (
    .a(\D1/LineCount [8]),
    .b(1'b0),
    .c(\D1/lt2_c8 ),
    .o({\D1/lt2_c9 ,open_n62}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt2_9  (
    .a(\D1/LineCount [9]),
    .b(1'b0),
    .c(\D1/lt2_c9 ),
    .o({\D1/lt2_c10 ,open_n63}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \D1/lt2_cin  (
    .a(1'b0),
    .o({\D1/lt2_c0 ,open_n66}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt2_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\D1/lt2_c16 ),
    .o({open_n67,LCD_SYNC_pad}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt3_0  (
    .a(\D1/PixelCount [0]),
    .b(1'b0),
    .c(\D1/lt3_c0 ),
    .o({\D1/lt3_c1 ,open_n68}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt3_1  (
    .a(\D1/PixelCount [1]),
    .b(1'b1),
    .c(\D1/lt3_c1 ),
    .o({\D1/lt3_c2 ,open_n69}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt3_10  (
    .a(\D1/PixelCount [10]),
    .b(1'b0),
    .c(\D1/lt3_c10 ),
    .o({\D1/lt3_c11 ,open_n70}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt3_11  (
    .a(\D1/PixelCount [11]),
    .b(1'b0),
    .c(\D1/lt3_c11 ),
    .o({\D1/lt3_c12 ,open_n71}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt3_12  (
    .a(\D1/PixelCount [12]),
    .b(1'b0),
    .c(\D1/lt3_c12 ),
    .o({\D1/lt3_c13 ,open_n72}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt3_13  (
    .a(\D1/PixelCount [13]),
    .b(1'b0),
    .c(\D1/lt3_c13 ),
    .o({\D1/lt3_c14 ,open_n73}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt3_14  (
    .a(\D1/PixelCount [14]),
    .b(1'b0),
    .c(\D1/lt3_c14 ),
    .o({\D1/lt3_c15 ,open_n74}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt3_15  (
    .a(\D1/PixelCount [15]),
    .b(1'b0),
    .c(\D1/lt3_c15 ),
    .o({\D1/lt3_c16 ,open_n75}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt3_2  (
    .a(\D1/PixelCount [2]),
    .b(1'b0),
    .c(\D1/lt3_c2 ),
    .o({\D1/lt3_c3 ,open_n76}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt3_3  (
    .a(\D1/PixelCount [3]),
    .b(1'b1),
    .c(\D1/lt3_c3 ),
    .o({\D1/lt3_c4 ,open_n77}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt3_4  (
    .a(\D1/PixelCount [4]),
    .b(1'b0),
    .c(\D1/lt3_c4 ),
    .o({\D1/lt3_c5 ,open_n78}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt3_5  (
    .a(\D1/PixelCount [5]),
    .b(1'b0),
    .c(\D1/lt3_c5 ),
    .o({\D1/lt3_c6 ,open_n79}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt3_6  (
    .a(\D1/PixelCount [6]),
    .b(1'b0),
    .c(\D1/lt3_c6 ),
    .o({\D1/lt3_c7 ,open_n80}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt3_7  (
    .a(\D1/PixelCount [7]),
    .b(1'b0),
    .c(\D1/lt3_c7 ),
    .o({\D1/lt3_c8 ,open_n81}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt3_8  (
    .a(\D1/PixelCount [8]),
    .b(1'b0),
    .c(\D1/lt3_c8 ),
    .o({\D1/lt3_c9 ,open_n82}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt3_9  (
    .a(\D1/PixelCount [9]),
    .b(1'b0),
    .c(\D1/lt3_c9 ),
    .o({\D1/lt3_c10 ,open_n83}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \D1/lt3_cin  (
    .a(1'b0),
    .o({\D1/lt3_c0 ,open_n86}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt3_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\D1/lt3_c16 ),
    .o({open_n87,FIFO_RST}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt4_0  (
    .a(1'b0),
    .b(\D1/PixelCount [0]),
    .c(\D1/lt4_c0 ),
    .o({\D1/lt4_c1 ,open_n88}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt4_1  (
    .a(1'b0),
    .b(\D1/PixelCount [1]),
    .c(\D1/lt4_c1 ),
    .o({\D1/lt4_c2 ,open_n89}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt4_10  (
    .a(1'b0),
    .b(\D1/PixelCount [10]),
    .c(\D1/lt4_c10 ),
    .o({\D1/lt4_c11 ,open_n90}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt4_11  (
    .a(1'b0),
    .b(\D1/PixelCount [11]),
    .c(\D1/lt4_c11 ),
    .o({\D1/lt4_c12 ,open_n91}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt4_12  (
    .a(1'b0),
    .b(\D1/PixelCount [12]),
    .c(\D1/lt4_c12 ),
    .o({\D1/lt4_c13 ,open_n92}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt4_13  (
    .a(1'b0),
    .b(\D1/PixelCount [13]),
    .c(\D1/lt4_c13 ),
    .o({\D1/lt4_c14 ,open_n93}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt4_14  (
    .a(1'b0),
    .b(\D1/PixelCount [14]),
    .c(\D1/lt4_c14 ),
    .o({\D1/lt4_c15 ,open_n94}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt4_15  (
    .a(1'b0),
    .b(\D1/PixelCount [15]),
    .c(\D1/lt4_c15 ),
    .o({\D1/lt4_c16 ,open_n95}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt4_2  (
    .a(1'b0),
    .b(\D1/PixelCount [2]),
    .c(\D1/lt4_c2 ),
    .o({\D1/lt4_c3 ,open_n96}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt4_3  (
    .a(1'b1),
    .b(\D1/PixelCount [3]),
    .c(\D1/lt4_c3 ),
    .o({\D1/lt4_c4 ,open_n97}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt4_4  (
    .a(1'b1),
    .b(\D1/PixelCount [4]),
    .c(\D1/lt4_c4 ),
    .o({\D1/lt4_c5 ,open_n98}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt4_5  (
    .a(1'b1),
    .b(\D1/PixelCount [5]),
    .c(\D1/lt4_c5 ),
    .o({\D1/lt4_c6 ,open_n99}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt4_6  (
    .a(1'b1),
    .b(\D1/PixelCount [6]),
    .c(\D1/lt4_c6 ),
    .o({\D1/lt4_c7 ,open_n100}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt4_7  (
    .a(1'b0),
    .b(\D1/PixelCount [7]),
    .c(\D1/lt4_c7 ),
    .o({\D1/lt4_c8 ,open_n101}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt4_8  (
    .a(1'b0),
    .b(\D1/PixelCount [8]),
    .c(\D1/lt4_c8 ),
    .o({\D1/lt4_c9 ,open_n102}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt4_9  (
    .a(1'b0),
    .b(\D1/PixelCount [9]),
    .c(\D1/lt4_c9 ),
    .o({\D1/lt4_c10 ,open_n103}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \D1/lt4_cin  (
    .a(1'b1),
    .o({\D1/lt4_c0 ,open_n106}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt4_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\D1/lt4_c16 ),
    .o({open_n107,\D1/n17 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt5_0  (
    .a(\D1/PixelCount [0]),
    .b(1'b0),
    .c(\D1/lt5_c0 ),
    .o({\D1/lt5_c1 ,open_n108}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt5_1  (
    .a(\D1/PixelCount [1]),
    .b(1'b0),
    .c(\D1/lt5_c1 ),
    .o({\D1/lt5_c2 ,open_n109}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt5_10  (
    .a(\D1/PixelCount [10]),
    .b(1'b0),
    .c(\D1/lt5_c10 ),
    .o({\D1/lt5_c11 ,open_n110}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt5_11  (
    .a(\D1/PixelCount [11]),
    .b(1'b0),
    .c(\D1/lt5_c11 ),
    .o({\D1/lt5_c12 ,open_n111}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt5_12  (
    .a(\D1/PixelCount [12]),
    .b(1'b0),
    .c(\D1/lt5_c12 ),
    .o({\D1/lt5_c13 ,open_n112}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt5_13  (
    .a(\D1/PixelCount [13]),
    .b(1'b0),
    .c(\D1/lt5_c13 ),
    .o({\D1/lt5_c14 ,open_n113}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt5_14  (
    .a(\D1/PixelCount [14]),
    .b(1'b0),
    .c(\D1/lt5_c14 ),
    .o({\D1/lt5_c15 ,open_n114}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt5_15  (
    .a(\D1/PixelCount [15]),
    .b(1'b0),
    .c(\D1/lt5_c15 ),
    .o({\D1/lt5_c16 ,open_n115}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt5_2  (
    .a(\D1/PixelCount [2]),
    .b(1'b0),
    .c(\D1/lt5_c2 ),
    .o({\D1/lt5_c3 ,open_n116}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt5_3  (
    .a(\D1/PixelCount [3]),
    .b(1'b0),
    .c(\D1/lt5_c3 ),
    .o({\D1/lt5_c4 ,open_n117}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt5_4  (
    .a(\D1/PixelCount [4]),
    .b(1'b1),
    .c(\D1/lt5_c4 ),
    .o({\D1/lt5_c5 ,open_n118}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt5_5  (
    .a(\D1/PixelCount [5]),
    .b(1'b0),
    .c(\D1/lt5_c5 ),
    .o({\D1/lt5_c6 ,open_n119}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt5_6  (
    .a(\D1/PixelCount [6]),
    .b(1'b1),
    .c(\D1/lt5_c6 ),
    .o({\D1/lt5_c7 ,open_n120}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt5_7  (
    .a(\D1/PixelCount [7]),
    .b(1'b1),
    .c(\D1/lt5_c7 ),
    .o({\D1/lt5_c8 ,open_n121}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt5_8  (
    .a(\D1/PixelCount [8]),
    .b(1'b0),
    .c(\D1/lt5_c8 ),
    .o({\D1/lt5_c9 ,open_n122}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt5_9  (
    .a(\D1/PixelCount [9]),
    .b(1'b1),
    .c(\D1/lt5_c9 ),
    .o({\D1/lt5_c10 ,open_n123}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \D1/lt5_cin  (
    .a(1'b1),
    .o({\D1/lt5_c0 ,open_n126}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt5_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\D1/lt5_c16 ),
    .o({open_n127,\D1/n18 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt6_0  (
    .a(1'b0),
    .b(\D1/LineCount [0]),
    .c(\D1/lt6_c0 ),
    .o({\D1/lt6_c1 ,open_n128}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt6_1  (
    .a(1'b1),
    .b(\D1/LineCount [1]),
    .c(\D1/lt6_c1 ),
    .o({\D1/lt6_c2 ,open_n129}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt6_10  (
    .a(1'b0),
    .b(\D1/LineCount [10]),
    .c(\D1/lt6_c10 ),
    .o({\D1/lt6_c11 ,open_n130}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt6_11  (
    .a(1'b0),
    .b(\D1/LineCount [11]),
    .c(\D1/lt6_c11 ),
    .o({\D1/lt6_c12 ,open_n131}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt6_12  (
    .a(1'b0),
    .b(\D1/LineCount [12]),
    .c(\D1/lt6_c12 ),
    .o({\D1/lt6_c13 ,open_n132}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt6_13  (
    .a(1'b0),
    .b(\D1/LineCount [13]),
    .c(\D1/lt6_c13 ),
    .o({\D1/lt6_c14 ,open_n133}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt6_14  (
    .a(1'b0),
    .b(\D1/LineCount [14]),
    .c(\D1/lt6_c14 ),
    .o({\D1/lt6_c15 ,open_n134}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt6_15  (
    .a(1'b0),
    .b(\D1/LineCount [15]),
    .c(\D1/lt6_c15 ),
    .o({\D1/lt6_c16 ,open_n135}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt6_2  (
    .a(1'b0),
    .b(\D1/LineCount [2]),
    .c(\D1/lt6_c2 ),
    .o({\D1/lt6_c3 ,open_n136}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt6_3  (
    .a(1'b1),
    .b(\D1/LineCount [3]),
    .c(\D1/lt6_c3 ),
    .o({\D1/lt6_c4 ,open_n137}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt6_4  (
    .a(1'b0),
    .b(\D1/LineCount [4]),
    .c(\D1/lt6_c4 ),
    .o({\D1/lt6_c5 ,open_n138}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt6_5  (
    .a(1'b0),
    .b(\D1/LineCount [5]),
    .c(\D1/lt6_c5 ),
    .o({\D1/lt6_c6 ,open_n139}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt6_6  (
    .a(1'b0),
    .b(\D1/LineCount [6]),
    .c(\D1/lt6_c6 ),
    .o({\D1/lt6_c7 ,open_n140}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt6_7  (
    .a(1'b0),
    .b(\D1/LineCount [7]),
    .c(\D1/lt6_c7 ),
    .o({\D1/lt6_c8 ,open_n141}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt6_8  (
    .a(1'b0),
    .b(\D1/LineCount [8]),
    .c(\D1/lt6_c8 ),
    .o({\D1/lt6_c9 ,open_n142}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt6_9  (
    .a(1'b0),
    .b(\D1/LineCount [9]),
    .c(\D1/lt6_c9 ),
    .o({\D1/lt6_c10 ,open_n143}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \D1/lt6_cin  (
    .a(1'b1),
    .o({\D1/lt6_c0 ,open_n146}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt6_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\D1/lt6_c16 ),
    .o({open_n147,\D1/n20 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt7_0  (
    .a(\D1/LineCount [0]),
    .b(1'b0),
    .c(\D1/lt7_c0 ),
    .o({\D1/lt7_c1 ,open_n148}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt7_1  (
    .a(\D1/LineCount [1]),
    .b(1'b0),
    .c(\D1/lt7_c1 ),
    .o({\D1/lt7_c2 ,open_n149}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt7_10  (
    .a(\D1/LineCount [10]),
    .b(1'b0),
    .c(\D1/lt7_c10 ),
    .o({\D1/lt7_c11 ,open_n150}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt7_11  (
    .a(\D1/LineCount [11]),
    .b(1'b0),
    .c(\D1/lt7_c11 ),
    .o({\D1/lt7_c12 ,open_n151}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt7_12  (
    .a(\D1/LineCount [12]),
    .b(1'b0),
    .c(\D1/lt7_c12 ),
    .o({\D1/lt7_c13 ,open_n152}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt7_13  (
    .a(\D1/LineCount [13]),
    .b(1'b0),
    .c(\D1/lt7_c13 ),
    .o({\D1/lt7_c14 ,open_n153}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt7_14  (
    .a(\D1/LineCount [14]),
    .b(1'b0),
    .c(\D1/lt7_c14 ),
    .o({\D1/lt7_c15 ,open_n154}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt7_15  (
    .a(\D1/LineCount [15]),
    .b(1'b0),
    .c(\D1/lt7_c15 ),
    .o({\D1/lt7_c16 ,open_n155}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt7_2  (
    .a(\D1/LineCount [2]),
    .b(1'b1),
    .c(\D1/lt7_c2 ),
    .o({\D1/lt7_c3 ,open_n156}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt7_3  (
    .a(\D1/LineCount [3]),
    .b(1'b0),
    .c(\D1/lt7_c3 ),
    .o({\D1/lt7_c4 ,open_n157}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt7_4  (
    .a(\D1/LineCount [4]),
    .b(1'b0),
    .c(\D1/lt7_c4 ),
    .o({\D1/lt7_c5 ,open_n158}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt7_5  (
    .a(\D1/LineCount [5]),
    .b(1'b1),
    .c(\D1/lt7_c5 ),
    .o({\D1/lt7_c6 ,open_n159}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt7_6  (
    .a(\D1/LineCount [6]),
    .b(1'b0),
    .c(\D1/lt7_c6 ),
    .o({\D1/lt7_c7 ,open_n160}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt7_7  (
    .a(\D1/LineCount [7]),
    .b(1'b0),
    .c(\D1/lt7_c7 ),
    .o({\D1/lt7_c8 ,open_n161}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt7_8  (
    .a(\D1/LineCount [8]),
    .b(1'b1),
    .c(\D1/lt7_c8 ),
    .o({\D1/lt7_c9 ,open_n162}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt7_9  (
    .a(\D1/LineCount [9]),
    .b(1'b0),
    .c(\D1/lt7_c9 ),
    .o({\D1/lt7_c10 ,open_n163}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \D1/lt7_cin  (
    .a(1'b0),
    .o({\D1/lt7_c0 ,open_n166}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt7_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\D1/lt7_c16 ),
    .o({open_n167,\D1/n22 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt8_0  (
    .a(1'b1),
    .b(\D1/PixelCount [0]),
    .c(\D1/lt8_c0 ),
    .o({\D1/lt8_c1 ,open_n168}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt8_1  (
    .a(1'b1),
    .b(\D1/PixelCount [1]),
    .c(\D1/lt8_c1 ),
    .o({\D1/lt8_c2 ,open_n169}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt8_10  (
    .a(1'b0),
    .b(\D1/PixelCount [10]),
    .c(\D1/lt8_c10 ),
    .o({\D1/lt8_c11 ,open_n170}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt8_11  (
    .a(1'b0),
    .b(\D1/PixelCount [11]),
    .c(\D1/lt8_c11 ),
    .o({\D1/lt8_c12 ,open_n171}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt8_12  (
    .a(1'b0),
    .b(\D1/PixelCount [12]),
    .c(\D1/lt8_c12 ),
    .o({\D1/lt8_c13 ,open_n172}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt8_13  (
    .a(1'b0),
    .b(\D1/PixelCount [13]),
    .c(\D1/lt8_c13 ),
    .o({\D1/lt8_c14 ,open_n173}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt8_14  (
    .a(1'b0),
    .b(\D1/PixelCount [14]),
    .c(\D1/lt8_c14 ),
    .o({\D1/lt8_c15 ,open_n174}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt8_15  (
    .a(1'b0),
    .b(\D1/PixelCount [15]),
    .c(\D1/lt8_c15 ),
    .o({\D1/lt8_c16 ,open_n175}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt8_2  (
    .a(1'b1),
    .b(\D1/PixelCount [2]),
    .c(\D1/lt8_c2 ),
    .o({\D1/lt8_c3 ,open_n176}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt8_3  (
    .a(1'b0),
    .b(\D1/PixelCount [3]),
    .c(\D1/lt8_c3 ),
    .o({\D1/lt8_c4 ,open_n177}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt8_4  (
    .a(1'b1),
    .b(\D1/PixelCount [4]),
    .c(\D1/lt8_c4 ),
    .o({\D1/lt8_c5 ,open_n178}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt8_5  (
    .a(1'b1),
    .b(\D1/PixelCount [5]),
    .c(\D1/lt8_c5 ),
    .o({\D1/lt8_c6 ,open_n179}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt8_6  (
    .a(1'b1),
    .b(\D1/PixelCount [6]),
    .c(\D1/lt8_c6 ),
    .o({\D1/lt8_c7 ,open_n180}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt8_7  (
    .a(1'b0),
    .b(\D1/PixelCount [7]),
    .c(\D1/lt8_c7 ),
    .o({\D1/lt8_c8 ,open_n181}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt8_8  (
    .a(1'b0),
    .b(\D1/PixelCount [8]),
    .c(\D1/lt8_c8 ),
    .o({\D1/lt8_c9 ,open_n182}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt8_9  (
    .a(1'b0),
    .b(\D1/PixelCount [9]),
    .c(\D1/lt8_c9 ),
    .o({\D1/lt8_c10 ,open_n183}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \D1/lt8_cin  (
    .a(1'b1),
    .o({\D1/lt8_c0 ,open_n186}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt8_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\D1/lt8_c16 ),
    .o({open_n187,\D1/n24 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt9_0  (
    .a(\D1/PixelCount [0]),
    .b(1'b1),
    .c(\D1/lt9_c0 ),
    .o({\D1/lt9_c1 ,open_n188}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt9_1  (
    .a(\D1/PixelCount [1]),
    .b(1'b0),
    .c(\D1/lt9_c1 ),
    .o({\D1/lt9_c2 ,open_n189}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt9_10  (
    .a(\D1/PixelCount [10]),
    .b(1'b0),
    .c(\D1/lt9_c10 ),
    .o({\D1/lt9_c11 ,open_n190}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt9_11  (
    .a(\D1/PixelCount [11]),
    .b(1'b0),
    .c(\D1/lt9_c11 ),
    .o({\D1/lt9_c12 ,open_n191}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt9_12  (
    .a(\D1/PixelCount [12]),
    .b(1'b0),
    .c(\D1/lt9_c12 ),
    .o({\D1/lt9_c13 ,open_n192}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt9_13  (
    .a(\D1/PixelCount [13]),
    .b(1'b0),
    .c(\D1/lt9_c13 ),
    .o({\D1/lt9_c14 ,open_n193}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt9_14  (
    .a(\D1/PixelCount [14]),
    .b(1'b0),
    .c(\D1/lt9_c14 ),
    .o({\D1/lt9_c15 ,open_n194}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt9_15  (
    .a(\D1/PixelCount [15]),
    .b(1'b0),
    .c(\D1/lt9_c15 ),
    .o({\D1/lt9_c16 ,open_n195}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt9_2  (
    .a(\D1/PixelCount [2]),
    .b(1'b0),
    .c(\D1/lt9_c2 ),
    .o({\D1/lt9_c3 ,open_n196}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt9_3  (
    .a(\D1/PixelCount [3]),
    .b(1'b1),
    .c(\D1/lt9_c3 ),
    .o({\D1/lt9_c4 ,open_n197}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt9_4  (
    .a(\D1/PixelCount [4]),
    .b(1'b1),
    .c(\D1/lt9_c4 ),
    .o({\D1/lt9_c5 ,open_n198}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt9_5  (
    .a(\D1/PixelCount [5]),
    .b(1'b0),
    .c(\D1/lt9_c5 ),
    .o({\D1/lt9_c6 ,open_n199}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt9_6  (
    .a(\D1/PixelCount [6]),
    .b(1'b1),
    .c(\D1/lt9_c6 ),
    .o({\D1/lt9_c7 ,open_n200}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt9_7  (
    .a(\D1/PixelCount [7]),
    .b(1'b0),
    .c(\D1/lt9_c7 ),
    .o({\D1/lt9_c8 ,open_n201}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt9_8  (
    .a(\D1/PixelCount [8]),
    .b(1'b0),
    .c(\D1/lt9_c8 ),
    .o({\D1/lt9_c9 ,open_n202}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt9_9  (
    .a(\D1/PixelCount [9]),
    .b(1'b1),
    .c(\D1/lt9_c9 ),
    .o({\D1/lt9_c10 ,open_n203}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \D1/lt9_cin  (
    .a(1'b1),
    .o({\D1/lt9_c0 ,open_n206}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \D1/lt9_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\D1/lt9_c16 ),
    .o({open_n207,\D1/n26 }));
  reg_ar_as_w1 \D1/reg0_b0  (
    .clk(LCD_CLK_pad),
    .d(\D1/n8 [0]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/PixelCount [0]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg0_b1  (
    .clk(LCD_CLK_pad),
    .d(\D1/n8 [1]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/PixelCount [1]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg0_b10  (
    .clk(LCD_CLK_pad),
    .d(\D1/n8 [10]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/PixelCount [10]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg0_b11  (
    .clk(LCD_CLK_pad),
    .d(\D1/n8 [11]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/PixelCount [11]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg0_b12  (
    .clk(LCD_CLK_pad),
    .d(\D1/n8 [12]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/PixelCount [12]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg0_b13  (
    .clk(LCD_CLK_pad),
    .d(\D1/n8 [13]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/PixelCount [13]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg0_b14  (
    .clk(LCD_CLK_pad),
    .d(\D1/n8 [14]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/PixelCount [14]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg0_b15  (
    .clk(LCD_CLK_pad),
    .d(\D1/n8 [15]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/PixelCount [15]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg0_b2  (
    .clk(LCD_CLK_pad),
    .d(\D1/n8 [2]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/PixelCount [2]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg0_b3  (
    .clk(LCD_CLK_pad),
    .d(\D1/n8 [3]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/PixelCount [3]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg0_b4  (
    .clk(LCD_CLK_pad),
    .d(\D1/n8 [4]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/PixelCount [4]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg0_b5  (
    .clk(LCD_CLK_pad),
    .d(\D1/n8 [5]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/PixelCount [5]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg0_b6  (
    .clk(LCD_CLK_pad),
    .d(\D1/n8 [6]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/PixelCount [6]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg0_b7  (
    .clk(LCD_CLK_pad),
    .d(\D1/n8 [7]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/PixelCount [7]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg0_b8  (
    .clk(LCD_CLK_pad),
    .d(\D1/n8 [8]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/PixelCount [8]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg0_b9  (
    .clk(LCD_CLK_pad),
    .d(\D1/n8 [9]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/PixelCount [9]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg1_b0  (
    .clk(LCD_CLK_pad),
    .d(\D1/n9 [0]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/LineCount [0]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg1_b1  (
    .clk(LCD_CLK_pad),
    .d(\D1/n9 [1]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/LineCount [1]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg1_b10  (
    .clk(LCD_CLK_pad),
    .d(\D1/n9 [10]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/LineCount [10]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg1_b11  (
    .clk(LCD_CLK_pad),
    .d(\D1/n9 [11]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/LineCount [11]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg1_b12  (
    .clk(LCD_CLK_pad),
    .d(\D1/n9 [12]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/LineCount [12]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg1_b13  (
    .clk(LCD_CLK_pad),
    .d(\D1/n9 [13]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/LineCount [13]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg1_b14  (
    .clk(LCD_CLK_pad),
    .d(\D1/n9 [14]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/LineCount [14]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg1_b15  (
    .clk(LCD_CLK_pad),
    .d(\D1/n9 [15]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/LineCount [15]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg1_b2  (
    .clk(LCD_CLK_pad),
    .d(\D1/n9 [2]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/LineCount [2]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg1_b3  (
    .clk(LCD_CLK_pad),
    .d(\D1/n9 [3]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/LineCount [3]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg1_b4  (
    .clk(LCD_CLK_pad),
    .d(\D1/n9 [4]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/LineCount [4]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg1_b5  (
    .clk(LCD_CLK_pad),
    .d(\D1/n9 [5]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/LineCount [5]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg1_b6  (
    .clk(LCD_CLK_pad),
    .d(\D1/n9 [6]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/LineCount [6]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg1_b7  (
    .clk(LCD_CLK_pad),
    .d(\D1/n9 [7]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/LineCount [7]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg1_b8  (
    .clk(LCD_CLK_pad),
    .d(\D1/n9 [8]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/LineCount [8]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  reg_ar_as_w1 \D1/reg1_b9  (
    .clk(LCD_CLK_pad),
    .d(\D1/n9 [9]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\D1/LineCount [9]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/VGAMod.v(72)
  EF2_PHY_FIFO #(
    .AE(32'b00000000000000000000000000110100),
    .AEP1(32'b00000000000000000000000000111100),
    .AF(32'b00000000000000000001111111101000),
    .AFM1(32'b00000000000000000001111111100100),
    .ASYNC_RESET_RELEASE("SYNC"),
    .DATA_WIDTH_A("4"),
    .DATA_WIDTH_B("9"),
    .E(32'b00000000000000000000000000000100),
    .EP1(32'b00000000000000000000000000001100),
    .F(32'b00000000000000000010000000000000),
    .FM1(32'b00000000000000000001111111111100),
    .GSR("DISABLE"),
    .MODE("FIFO8K"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"))
    \FIFO0/logic_fifo_0  (
    .clkr(LCD_CLK_pad),
    .clkw(FIFO_CLK_W),
    .csr({2'b11,\D1/n28 }),
    .csw({2'b11,\FIFO0/logic_fifo_full_neg }),
    .dia({open_n208,open_n209,open_n210,open_n211,open_n212,FIFO_DI[3:0]}),
    .orea(1'b0),
    .oreb(1'b0),
    .re(FIFO_RE),
    .rprst(FIFO_RST),
    .rst(FIFO_RST),
    .we(FIFO_WE),
    .dob({open_n233,FIFO_DO[3:0],FIFO_DO[11:8]}),
    .empty_flag(FIFO_EMPTY),
    .full_flag(\FIFO0/logic_fifo_full ));
  EF2_PHY_FIFO #(
    .AE(32'b00000000000000000000000000110100),
    .AEP1(32'b00000000000000000000000000111100),
    .AF(32'b00000000000000000001111111101000),
    .AFM1(32'b00000000000000000001111111100100),
    .ASYNC_RESET_RELEASE("SYNC"),
    .DATA_WIDTH_A("4"),
    .DATA_WIDTH_B("9"),
    .E(32'b00000000000000000000000000000100),
    .EP1(32'b00000000000000000000000000001100),
    .F(32'b00000000000000000010000000000000),
    .FM1(32'b00000000000000000001111111111100),
    .GSR("DISABLE"),
    .MODE("FIFO8K"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("ASYNC"))
    \FIFO0/logic_fifo_1  (
    .clkr(LCD_CLK_pad),
    .clkw(FIFO_CLK_W),
    .csr({2'b11,\D1/n28 }),
    .csw({2'b11,\FIFO0/logic_fifo_full_neg }),
    .dia({open_n234,open_n235,open_n236,open_n237,open_n238,FIFO_DI[7:4]}),
    .orea(1'b0),
    .oreb(1'b0),
    .re(FIFO_RE),
    .rprst(FIFO_RST),
    .rst(FIFO_RST),
    .we(FIFO_WE),
    .dob({open_n259,FIFO_DO[7:4],FIFO_DO[15:12]}));
  EF2_PHY_GCLK \PLL1/bufg_feedback  (
    .clki(\PLL1/clk0_buf ),
    .clko(CLK_100M));  // al_ip/LCDPLL.v(41)
  EF2_PHY_PLL #(
    .CLKC0_CPHASE(9),
    .CLKC0_DIV(10),
    .CLKC0_DIV2_ENABLE("DISABLE"),
    .CLKC0_DUTY(0.500000),
    .CLKC0_DUTY50("ENABLE"),
    .CLKC0_DUTY_INT(5),
    .CLKC0_ENABLE("ENABLE"),
    .CLKC0_FPHASE(0),
    .CLKC1_CPHASE(29),
    .CLKC1_DIV(30),
    .CLKC1_DIV2_ENABLE("DISABLE"),
    .CLKC1_DUTY(0.500000),
    .CLKC1_DUTY50("ENABLE"),
    .CLKC1_DUTY_INT(15),
    .CLKC1_ENABLE("ENABLE"),
    .CLKC1_FPHASE(0),
    .CLKC2_CPHASE(39),
    .CLKC2_DIV(40),
    .CLKC2_DIV2_ENABLE("DISABLE"),
    .CLKC2_ENABLE("ENABLE"),
    .CLKC2_FPHASE(0),
    .CLKC3_CPHASE(110),
    .CLKC3_DIV(111),
    .CLKC3_DIV2_ENABLE("DISABLE"),
    .CLKC3_ENABLE("ENABLE"),
    .CLKC3_FPHASE(0),
    .CLKC4_CPHASE(1),
    .CLKC4_DIV(1),
    .CLKC4_DIV2_ENABLE("DISABLE"),
    .CLKC4_ENABLE("DISABLE"),
    .CLKC4_FPHASE(0),
    .CLKC5_CPHASE(1),
    .CLKC5_DIV(1),
    .CLKC5_DIV2_ENABLE("DISABLE"),
    .CLKC5_ENABLE("DISABLE"),
    .CLKC6_CPHASE(1),
    .CLKC6_DIV(1),
    .CLKC6_DIV2_ENABLE("DISABLE"),
    .CLKC6_ENABLE("DISABLE"),
    .DERIVE_PLL_CLOCKS("DISABLE"),
    .DPHASE_SOURCE("DISABLE"),
    .DYNCFG("DISABLE"),
    .FBCLK_DIV(6),
    .FEEDBK_MODE("NORMAL"),
    .FEEDBK_PATH("CLKC0_EXT"),
    .FIN("50.000"),
    .FREQ_LOCK_ACCURACY(2),
    .FREQ_OFFSET("0.000000"),
    .FREQ_OFFSET_INT("0"),
    .GEN_BASIC_CLOCK("DISABLE"),
    .GMC_GAIN(6),
    .GMC_TEST(14),
    .HIGH_SPEED_EN("ENABLE"),
    .ICP_CURRENT(3),
    .IF_ESCLKSTSW("DISABLE"),
    .INTFB_WAKE("DISABLE"),
    .INTPI(3),
    .KVCO(6),
    .LPF_CAPACITOR(3),
    .LPF_RESISTOR(2),
    .NORESET("DISABLE"),
    .ODIV_MUXC0("DIV"),
    .ODIV_MUXC1("DIV"),
    .ODIV_MUXC2("DIV"),
    .ODIV_MUXC3("DIV"),
    .ODIV_MUXC4("DIV"),
    .OFFSET_MODE("EXT"),
    .PLLC2RST_ENA("DISABLE"),
    .PLLC34RST_ENA("DISABLE"),
    .PLLMRST_ENA("DISABLE"),
    .PLLRST_ENA("ENABLE"),
    .PLL_LOCK_MODE(0),
    .PREDIV_MUXC0("VCO"),
    .PREDIV_MUXC1("VCO"),
    .PREDIV_MUXC2("VCO"),
    .PREDIV_MUXC3("VCO"),
    .PREDIV_MUXC4("VCO"),
    .PREDIV_MUXC5("VCO"),
    .PREDIV_MUXC6("VCO"),
    .PU_INTP("DISABLE"),
    .REFCLK_DIV(3),
    .REFCLK_SEL("INTERNAL"),
    .SSC_AMP("0.000000"),
    .SSC_ENABLE("DISABLE"),
    .SSC_FREQ_DIV(0),
    .SSC_MODE("Down"),
    .SSC_RNGE(0),
    .STDBY_ENABLE("DISABLE"),
    .STDBY_VCO_ENA("DISABLE"),
    .SYNC_ENABLE("DISABLE"),
    .VCO_NORESET("DISABLE"))
    \PLL1/pll_inst  (
    .daddr(6'b000000),
    .dclk(1'b0),
    .dcs(1'b0),
    .di(8'b00000000),
    .dsm_refclk(1'b0),
    .dsm_rst(1'b0),
    .dwe(1'b0),
    .fbclk(CLK_100M),
    .frac_offset_valid(1'b0),
    .psclk(1'b0),
    .psclksel(3'b000),
    .psdown(1'b0),
    .psstep(1'b0),
    .refclk(clk_pad),
    .reset(1'b0),
    .ssc_en(1'b0),
    .stdby(1'b0),
    .clkc({open_n262,open_n263,open_n264,LCD_CLK_pad,open_n265,open_n266,\PLL1/clk0_buf }));  // al_ip/LCDPLL.v(93)
  reg_ar_as_w1 \U1/CLK_OUT_reg  (
    .clk(LCD_CLK_pad),
    .d(\U1/n2 ),
    .en(\U1/n1 ),
    .reset(1'b0),
    .set(~nRST_pad),
    .q(LED_pad[0]));  // source/CLK_MOD.v(32)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u0  (
    .a(\U1/Count [0]),
    .b(1'b1),
    .c(\U1/add0/c0 ),
    .o({\U1/add0/c1 ,\U1/n3 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u1  (
    .a(\U1/Count [1]),
    .b(1'b0),
    .c(\U1/add0/c1 ),
    .o({\U1/add0/c2 ,\U1/n3 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u10  (
    .a(\U1/Count [10]),
    .b(1'b0),
    .c(\U1/add0/c10 ),
    .o({\U1/add0/c11 ,\U1/n3 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u11  (
    .a(\U1/Count [11]),
    .b(1'b0),
    .c(\U1/add0/c11 ),
    .o({\U1/add0/c12 ,\U1/n3 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u12  (
    .a(\U1/Count [12]),
    .b(1'b0),
    .c(\U1/add0/c12 ),
    .o({\U1/add0/c13 ,\U1/n3 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u13  (
    .a(\U1/Count [13]),
    .b(1'b0),
    .c(\U1/add0/c13 ),
    .o({\U1/add0/c14 ,\U1/n3 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u14  (
    .a(\U1/Count [14]),
    .b(1'b0),
    .c(\U1/add0/c14 ),
    .o({\U1/add0/c15 ,\U1/n3 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u15  (
    .a(\U1/Count [15]),
    .b(1'b0),
    .c(\U1/add0/c15 ),
    .o({\U1/add0/c16 ,\U1/n3 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u16  (
    .a(\U1/Count [16]),
    .b(1'b0),
    .c(\U1/add0/c16 ),
    .o({\U1/add0/c17 ,\U1/n3 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u17  (
    .a(\U1/Count [17]),
    .b(1'b0),
    .c(\U1/add0/c17 ),
    .o({\U1/add0/c18 ,\U1/n3 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u18  (
    .a(\U1/Count [18]),
    .b(1'b0),
    .c(\U1/add0/c18 ),
    .o({\U1/add0/c19 ,\U1/n3 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u19  (
    .a(\U1/Count [19]),
    .b(1'b0),
    .c(\U1/add0/c19 ),
    .o({\U1/add0/c20 ,\U1/n3 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u2  (
    .a(\U1/Count [2]),
    .b(1'b0),
    .c(\U1/add0/c2 ),
    .o({\U1/add0/c3 ,\U1/n3 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u20  (
    .a(\U1/Count [20]),
    .b(1'b0),
    .c(\U1/add0/c20 ),
    .o({\U1/add0/c21 ,\U1/n3 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u21  (
    .a(\U1/Count [21]),
    .b(1'b0),
    .c(\U1/add0/c21 ),
    .o({\U1/add0/c22 ,\U1/n3 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u22  (
    .a(\U1/Count [22]),
    .b(1'b0),
    .c(\U1/add0/c22 ),
    .o({\U1/add0/c23 ,\U1/n3 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u23  (
    .a(\U1/Count [23]),
    .b(1'b0),
    .c(\U1/add0/c23 ),
    .o({\U1/add0/c24 ,\U1/n3 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u24  (
    .a(\U1/Count [24]),
    .b(1'b0),
    .c(\U1/add0/c24 ),
    .o({\U1/add0/c25 ,\U1/n3 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u25  (
    .a(\U1/Count [25]),
    .b(1'b0),
    .c(\U1/add0/c25 ),
    .o({\U1/add0/c26 ,\U1/n3 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u26  (
    .a(\U1/Count [26]),
    .b(1'b0),
    .c(\U1/add0/c26 ),
    .o({\U1/add0/c27 ,\U1/n3 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u27  (
    .a(\U1/Count [27]),
    .b(1'b0),
    .c(\U1/add0/c27 ),
    .o({\U1/add0/c28 ,\U1/n3 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u28  (
    .a(\U1/Count [28]),
    .b(1'b0),
    .c(\U1/add0/c28 ),
    .o({\U1/add0/c29 ,\U1/n3 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u29  (
    .a(\U1/Count [29]),
    .b(1'b0),
    .c(\U1/add0/c29 ),
    .o({\U1/add0/c30 ,\U1/n3 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u3  (
    .a(\U1/Count [3]),
    .b(1'b0),
    .c(\U1/add0/c3 ),
    .o({\U1/add0/c4 ,\U1/n3 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u30  (
    .a(\U1/Count [30]),
    .b(1'b0),
    .c(\U1/add0/c30 ),
    .o({\U1/add0/c31 ,\U1/n3 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u31  (
    .a(\U1/Count [31]),
    .b(1'b0),
    .c(\U1/add0/c31 ),
    .o({open_n277,\U1/n3 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u4  (
    .a(\U1/Count [4]),
    .b(1'b0),
    .c(\U1/add0/c4 ),
    .o({\U1/add0/c5 ,\U1/n3 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u5  (
    .a(\U1/Count [5]),
    .b(1'b0),
    .c(\U1/add0/c5 ),
    .o({\U1/add0/c6 ,\U1/n3 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u6  (
    .a(\U1/Count [6]),
    .b(1'b0),
    .c(\U1/add0/c6 ),
    .o({\U1/add0/c7 ,\U1/n3 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u7  (
    .a(\U1/Count [7]),
    .b(1'b0),
    .c(\U1/add0/c7 ),
    .o({\U1/add0/c8 ,\U1/n3 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u8  (
    .a(\U1/Count [8]),
    .b(1'b0),
    .c(\U1/add0/c8 ),
    .o({\U1/add0/c9 ,\U1/n3 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U1/add0/u9  (
    .a(\U1/Count [9]),
    .b(1'b0),
    .c(\U1/add0/c9 ),
    .o({\U1/add0/c10 ,\U1/n3 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \U1/add0/ucin  (
    .a(1'b0),
    .o({\U1/add0/c0 ,open_n280}));
  reg_ar_as_w1 \U1/reg0_b0  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [0]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [0]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b1  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [1]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [1]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b10  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [10]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [10]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b11  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [11]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [11]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b12  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [12]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [12]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b13  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [13]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [13]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b14  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [14]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [14]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b15  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [15]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [15]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b16  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [16]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [16]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b17  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [17]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [17]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b18  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [18]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [18]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b19  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [19]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [19]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b2  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [2]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [2]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b20  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [20]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [20]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b21  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [21]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [21]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b22  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [22]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [22]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b23  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [23]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [23]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b24  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [24]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [24]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b25  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [25]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [25]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b26  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [26]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [26]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b27  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [27]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [27]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b28  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [28]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [28]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b29  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [29]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [29]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b3  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [3]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [3]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b30  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [30]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [30]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b31  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [31]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [31]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b4  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [4]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [4]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b5  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [5]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [5]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b6  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [6]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [6]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b7  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [7]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [7]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b8  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [8]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [8]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U1/reg0_b9  (
    .clk(LCD_CLK_pad),
    .d(\U1/n5 [9]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U1/Count [9]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/CLK_OUT_reg  (
    .clk(clk_pad),
    .d(\U2/n2 ),
    .en(\U2/n1 ),
    .reset(1'b0),
    .set(~nRST_pad),
    .q(LED_pad[1]));  // source/CLK_MOD.v(32)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u0  (
    .a(\U2/Count [0]),
    .b(1'b1),
    .c(\U2/add0/c0 ),
    .o({\U2/add0/c1 ,\U2/n3 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u1  (
    .a(\U2/Count [1]),
    .b(1'b0),
    .c(\U2/add0/c1 ),
    .o({\U2/add0/c2 ,\U2/n3 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u10  (
    .a(\U2/Count [10]),
    .b(1'b0),
    .c(\U2/add0/c10 ),
    .o({\U2/add0/c11 ,\U2/n3 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u11  (
    .a(\U2/Count [11]),
    .b(1'b0),
    .c(\U2/add0/c11 ),
    .o({\U2/add0/c12 ,\U2/n3 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u12  (
    .a(\U2/Count [12]),
    .b(1'b0),
    .c(\U2/add0/c12 ),
    .o({\U2/add0/c13 ,\U2/n3 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u13  (
    .a(\U2/Count [13]),
    .b(1'b0),
    .c(\U2/add0/c13 ),
    .o({\U2/add0/c14 ,\U2/n3 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u14  (
    .a(\U2/Count [14]),
    .b(1'b0),
    .c(\U2/add0/c14 ),
    .o({\U2/add0/c15 ,\U2/n3 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u15  (
    .a(\U2/Count [15]),
    .b(1'b0),
    .c(\U2/add0/c15 ),
    .o({\U2/add0/c16 ,\U2/n3 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u16  (
    .a(\U2/Count [16]),
    .b(1'b0),
    .c(\U2/add0/c16 ),
    .o({\U2/add0/c17 ,\U2/n3 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u17  (
    .a(\U2/Count [17]),
    .b(1'b0),
    .c(\U2/add0/c17 ),
    .o({\U2/add0/c18 ,\U2/n3 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u18  (
    .a(\U2/Count [18]),
    .b(1'b0),
    .c(\U2/add0/c18 ),
    .o({\U2/add0/c19 ,\U2/n3 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u19  (
    .a(\U2/Count [19]),
    .b(1'b0),
    .c(\U2/add0/c19 ),
    .o({\U2/add0/c20 ,\U2/n3 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u2  (
    .a(\U2/Count [2]),
    .b(1'b0),
    .c(\U2/add0/c2 ),
    .o({\U2/add0/c3 ,\U2/n3 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u20  (
    .a(\U2/Count [20]),
    .b(1'b0),
    .c(\U2/add0/c20 ),
    .o({\U2/add0/c21 ,\U2/n3 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u21  (
    .a(\U2/Count [21]),
    .b(1'b0),
    .c(\U2/add0/c21 ),
    .o({\U2/add0/c22 ,\U2/n3 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u22  (
    .a(\U2/Count [22]),
    .b(1'b0),
    .c(\U2/add0/c22 ),
    .o({\U2/add0/c23 ,\U2/n3 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u23  (
    .a(\U2/Count [23]),
    .b(1'b0),
    .c(\U2/add0/c23 ),
    .o({\U2/add0/c24 ,\U2/n3 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u24  (
    .a(\U2/Count [24]),
    .b(1'b0),
    .c(\U2/add0/c24 ),
    .o({\U2/add0/c25 ,\U2/n3 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u25  (
    .a(\U2/Count [25]),
    .b(1'b0),
    .c(\U2/add0/c25 ),
    .o({\U2/add0/c26 ,\U2/n3 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u26  (
    .a(\U2/Count [26]),
    .b(1'b0),
    .c(\U2/add0/c26 ),
    .o({\U2/add0/c27 ,\U2/n3 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u27  (
    .a(\U2/Count [27]),
    .b(1'b0),
    .c(\U2/add0/c27 ),
    .o({\U2/add0/c28 ,\U2/n3 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u28  (
    .a(\U2/Count [28]),
    .b(1'b0),
    .c(\U2/add0/c28 ),
    .o({\U2/add0/c29 ,\U2/n3 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u29  (
    .a(\U2/Count [29]),
    .b(1'b0),
    .c(\U2/add0/c29 ),
    .o({\U2/add0/c30 ,\U2/n3 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u3  (
    .a(\U2/Count [3]),
    .b(1'b0),
    .c(\U2/add0/c3 ),
    .o({\U2/add0/c4 ,\U2/n3 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u30  (
    .a(\U2/Count [30]),
    .b(1'b0),
    .c(\U2/add0/c30 ),
    .o({\U2/add0/c31 ,\U2/n3 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u31  (
    .a(\U2/Count [31]),
    .b(1'b0),
    .c(\U2/add0/c31 ),
    .o({open_n281,\U2/n3 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u4  (
    .a(\U2/Count [4]),
    .b(1'b0),
    .c(\U2/add0/c4 ),
    .o({\U2/add0/c5 ,\U2/n3 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u5  (
    .a(\U2/Count [5]),
    .b(1'b0),
    .c(\U2/add0/c5 ),
    .o({\U2/add0/c6 ,\U2/n3 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u6  (
    .a(\U2/Count [6]),
    .b(1'b0),
    .c(\U2/add0/c6 ),
    .o({\U2/add0/c7 ,\U2/n3 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u7  (
    .a(\U2/Count [7]),
    .b(1'b0),
    .c(\U2/add0/c7 ),
    .o({\U2/add0/c8 ,\U2/n3 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u8  (
    .a(\U2/Count [8]),
    .b(1'b0),
    .c(\U2/add0/c8 ),
    .o({\U2/add0/c9 ,\U2/n3 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U2/add0/u9  (
    .a(\U2/Count [9]),
    .b(1'b0),
    .c(\U2/add0/c9 ),
    .o({\U2/add0/c10 ,\U2/n3 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \U2/add0/ucin  (
    .a(1'b0),
    .o({\U2/add0/c0 ,open_n284}));
  reg_ar_as_w1 \U2/reg0_b0  (
    .clk(clk_pad),
    .d(\U2/n5 [0]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [0]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b1  (
    .clk(clk_pad),
    .d(\U2/n5 [1]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [1]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b10  (
    .clk(clk_pad),
    .d(\U2/n5 [10]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [10]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b11  (
    .clk(clk_pad),
    .d(\U2/n5 [11]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [11]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b12  (
    .clk(clk_pad),
    .d(\U2/n5 [12]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [12]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b13  (
    .clk(clk_pad),
    .d(\U2/n5 [13]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [13]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b14  (
    .clk(clk_pad),
    .d(\U2/n5 [14]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [14]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b15  (
    .clk(clk_pad),
    .d(\U2/n5 [15]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [15]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b16  (
    .clk(clk_pad),
    .d(\U2/n5 [16]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [16]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b17  (
    .clk(clk_pad),
    .d(\U2/n5 [17]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [17]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b18  (
    .clk(clk_pad),
    .d(\U2/n5 [18]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [18]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b19  (
    .clk(clk_pad),
    .d(\U2/n5 [19]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [19]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b2  (
    .clk(clk_pad),
    .d(\U2/n5 [2]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [2]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b20  (
    .clk(clk_pad),
    .d(\U2/n5 [20]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [20]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b21  (
    .clk(clk_pad),
    .d(\U2/n5 [21]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [21]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b22  (
    .clk(clk_pad),
    .d(\U2/n5 [22]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [22]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b23  (
    .clk(clk_pad),
    .d(\U2/n5 [23]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [23]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b24  (
    .clk(clk_pad),
    .d(\U2/n5 [24]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [24]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b25  (
    .clk(clk_pad),
    .d(\U2/n5 [25]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [25]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b26  (
    .clk(clk_pad),
    .d(\U2/n5 [26]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [26]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b27  (
    .clk(clk_pad),
    .d(\U2/n5 [27]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [27]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b28  (
    .clk(clk_pad),
    .d(\U2/n5 [28]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [28]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b29  (
    .clk(clk_pad),
    .d(\U2/n5 [29]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [29]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b3  (
    .clk(clk_pad),
    .d(\U2/n5 [3]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [3]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b30  (
    .clk(clk_pad),
    .d(\U2/n5 [30]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [30]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b31  (
    .clk(clk_pad),
    .d(\U2/n5 [31]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [31]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b4  (
    .clk(clk_pad),
    .d(\U2/n5 [4]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [4]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b5  (
    .clk(clk_pad),
    .d(\U2/n5 [5]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [5]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b6  (
    .clk(clk_pad),
    .d(\U2/n5 [6]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [6]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b7  (
    .clk(clk_pad),
    .d(\U2/n5 [7]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [7]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b8  (
    .clk(clk_pad),
    .d(\U2/n5 [8]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [8]));  // source/CLK_MOD.v(32)
  reg_ar_as_w1 \U2/reg0_b9  (
    .clk(clk_pad),
    .d(\U2/n5 [9]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U2/Count [9]));  // source/CLK_MOD.v(32)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U4/add0/u0  (
    .a(\U4/AddrCtrl [0]),
    .b(1'b1),
    .c(\U4/add0/c0 ),
    .o({\U4/add0/c1 ,\U4/n18 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U4/add0/u1  (
    .a(\U4/AddrCtrl [1]),
    .b(1'b0),
    .c(\U4/add0/c1 ),
    .o({\U4/add0/c2 ,\U4/n18 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U4/add0/u10  (
    .a(\U4/AddrCtrl [10]),
    .b(1'b0),
    .c(\U4/add0/c10 ),
    .o({\U4/add0/c11 ,\U4/n18 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U4/add0/u11  (
    .a(\U4/AddrCtrl [11]),
    .b(1'b0),
    .c(\U4/add0/c11 ),
    .o({\U4/add0/c12 ,\U4/n18 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U4/add0/u12  (
    .a(\U4/AddrCtrl [12]),
    .b(1'b0),
    .c(\U4/add0/c12 ),
    .o({\U4/add0/c13 ,\U4/n18 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U4/add0/u13  (
    .a(\U4/AddrCtrl [13]),
    .b(1'b0),
    .c(\U4/add0/c13 ),
    .o({\U4/add0/c14 ,\U4/n18 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U4/add0/u14  (
    .a(\U4/AddrCtrl [14]),
    .b(1'b0),
    .c(\U4/add0/c14 ),
    .o({\U4/add0/c15 ,\U4/n18 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U4/add0/u15  (
    .a(\U4/AddrCtrl [15]),
    .b(1'b0),
    .c(\U4/add0/c15 ),
    .o({open_n285,\U4/n18 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U4/add0/u2  (
    .a(\U4/AddrCtrl [2]),
    .b(1'b0),
    .c(\U4/add0/c2 ),
    .o({\U4/add0/c3 ,\U4/n18 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U4/add0/u3  (
    .a(\U4/AddrCtrl [3]),
    .b(1'b0),
    .c(\U4/add0/c3 ),
    .o({\U4/add0/c4 ,\U4/n18 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U4/add0/u4  (
    .a(\U4/AddrCtrl [4]),
    .b(1'b0),
    .c(\U4/add0/c4 ),
    .o({\U4/add0/c5 ,\U4/n18 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U4/add0/u5  (
    .a(\U4/AddrCtrl [5]),
    .b(1'b0),
    .c(\U4/add0/c5 ),
    .o({\U4/add0/c6 ,\U4/n18 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U4/add0/u6  (
    .a(\U4/AddrCtrl [6]),
    .b(1'b0),
    .c(\U4/add0/c6 ),
    .o({\U4/add0/c7 ,\U4/n18 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U4/add0/u7  (
    .a(\U4/AddrCtrl [7]),
    .b(1'b0),
    .c(\U4/add0/c7 ),
    .o({\U4/add0/c8 ,\U4/n18 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U4/add0/u8  (
    .a(\U4/AddrCtrl [8]),
    .b(1'b0),
    .c(\U4/add0/c8 ),
    .o({\U4/add0/c9 ,\U4/n18 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \U4/add0/u9  (
    .a(\U4/AddrCtrl [9]),
    .b(1'b0),
    .c(\U4/add0/c9 ),
    .o({\U4/add0/c10 ,\U4/n18 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \U4/add0/ucin  (
    .a(1'b0),
    .o({\U4/add0/c0 ,open_n288}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt0_0  (
    .a(\U4/AddrCtrl [0]),
    .b(1'b0),
    .c(\U4/lt0_c0 ),
    .o({\U4/lt0_c1 ,open_n289}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt0_1  (
    .a(\U4/AddrCtrl [1]),
    .b(1'b0),
    .c(\U4/lt0_c1 ),
    .o({\U4/lt0_c2 ,open_n290}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt0_10  (
    .a(\U4/AddrCtrl [10]),
    .b(1'b1),
    .c(\U4/lt0_c10 ),
    .o({\U4/lt0_c11 ,open_n291}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt0_11  (
    .a(\U4/AddrCtrl [11]),
    .b(1'b0),
    .c(\U4/lt0_c11 ),
    .o({\U4/lt0_c12 ,open_n292}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt0_12  (
    .a(\U4/AddrCtrl [12]),
    .b(1'b0),
    .c(\U4/lt0_c12 ),
    .o({\U4/lt0_c13 ,open_n293}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt0_13  (
    .a(\U4/AddrCtrl [13]),
    .b(1'b0),
    .c(\U4/lt0_c13 ),
    .o({\U4/lt0_c14 ,open_n294}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt0_14  (
    .a(\U4/AddrCtrl [14]),
    .b(1'b0),
    .c(\U4/lt0_c14 ),
    .o({\U4/lt0_c15 ,open_n295}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt0_15  (
    .a(\U4/AddrCtrl [15]),
    .b(1'b0),
    .c(\U4/lt0_c15 ),
    .o({\U4/lt0_c16 ,open_n296}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt0_2  (
    .a(\U4/AddrCtrl [2]),
    .b(1'b0),
    .c(\U4/lt0_c2 ),
    .o({\U4/lt0_c3 ,open_n297}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt0_3  (
    .a(\U4/AddrCtrl [3]),
    .b(1'b0),
    .c(\U4/lt0_c3 ),
    .o({\U4/lt0_c4 ,open_n298}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt0_4  (
    .a(\U4/AddrCtrl [4]),
    .b(1'b1),
    .c(\U4/lt0_c4 ),
    .o({\U4/lt0_c5 ,open_n299}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt0_5  (
    .a(\U4/AddrCtrl [5]),
    .b(1'b0),
    .c(\U4/lt0_c5 ),
    .o({\U4/lt0_c6 ,open_n300}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt0_6  (
    .a(\U4/AddrCtrl [6]),
    .b(1'b1),
    .c(\U4/lt0_c6 ),
    .o({\U4/lt0_c7 ,open_n301}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt0_7  (
    .a(\U4/AddrCtrl [7]),
    .b(1'b1),
    .c(\U4/lt0_c7 ),
    .o({\U4/lt0_c8 ,open_n302}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt0_8  (
    .a(\U4/AddrCtrl [8]),
    .b(1'b1),
    .c(\U4/lt0_c8 ),
    .o({\U4/lt0_c9 ,open_n303}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt0_9  (
    .a(\U4/AddrCtrl [9]),
    .b(1'b1),
    .c(\U4/lt0_c9 ),
    .o({\U4/lt0_c10 ,open_n304}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \U4/lt0_cin  (
    .a(1'b0),
    .o({\U4/lt0_c0 ,open_n307}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt0_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\U4/lt0_c16 ),
    .o({open_n308,\U4/n17 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt1_0  (
    .a(\U4/AddrCtrl [0]),
    .b(1'b0),
    .c(\U4/lt1_c0 ),
    .o({\U4/lt1_c1 ,open_n309}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt1_1  (
    .a(\U4/AddrCtrl [1]),
    .b(1'b0),
    .c(\U4/lt1_c1 ),
    .o({\U4/lt1_c2 ,open_n310}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt1_10  (
    .a(\U4/AddrCtrl [10]),
    .b(1'b1),
    .c(\U4/lt1_c10 ),
    .o({\U4/lt1_c11 ,open_n311}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt1_11  (
    .a(\U4/AddrCtrl [11]),
    .b(1'b0),
    .c(\U4/lt1_c11 ),
    .o({\U4/lt1_c12 ,open_n312}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt1_12  (
    .a(\U4/AddrCtrl [12]),
    .b(1'b0),
    .c(\U4/lt1_c12 ),
    .o({\U4/lt1_c13 ,open_n313}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt1_13  (
    .a(\U4/AddrCtrl [13]),
    .b(1'b0),
    .c(\U4/lt1_c13 ),
    .o({\U4/lt1_c14 ,open_n314}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt1_14  (
    .a(\U4/AddrCtrl [14]),
    .b(1'b0),
    .c(\U4/lt1_c14 ),
    .o({\U4/lt1_c15 ,open_n315}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt1_15  (
    .a(\U4/AddrCtrl [15]),
    .b(1'b0),
    .c(\U4/lt1_c15 ),
    .o({\U4/lt1_c16 ,open_n316}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt1_2  (
    .a(\U4/AddrCtrl [2]),
    .b(1'b0),
    .c(\U4/lt1_c2 ),
    .o({\U4/lt1_c3 ,open_n317}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt1_3  (
    .a(\U4/AddrCtrl [3]),
    .b(1'b0),
    .c(\U4/lt1_c3 ),
    .o({\U4/lt1_c4 ,open_n318}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt1_4  (
    .a(\U4/AddrCtrl [4]),
    .b(1'b0),
    .c(\U4/lt1_c4 ),
    .o({\U4/lt1_c5 ,open_n319}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt1_5  (
    .a(\U4/AddrCtrl [5]),
    .b(1'b0),
    .c(\U4/lt1_c5 ),
    .o({\U4/lt1_c6 ,open_n320}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt1_6  (
    .a(\U4/AddrCtrl [6]),
    .b(1'b1),
    .c(\U4/lt1_c6 ),
    .o({\U4/lt1_c7 ,open_n321}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt1_7  (
    .a(\U4/AddrCtrl [7]),
    .b(1'b0),
    .c(\U4/lt1_c7 ),
    .o({\U4/lt1_c8 ,open_n322}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt1_8  (
    .a(\U4/AddrCtrl [8]),
    .b(1'b0),
    .c(\U4/lt1_c8 ),
    .o({\U4/lt1_c9 ,open_n323}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt1_9  (
    .a(\U4/AddrCtrl [9]),
    .b(1'b1),
    .c(\U4/lt1_c9 ),
    .o({\U4/lt1_c10 ,open_n324}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \U4/lt1_cin  (
    .a(1'b0),
    .o({\U4/lt1_c0 ,open_n327}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt1_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\U4/lt1_c16 ),
    .o({open_n328,\U4/n23 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt2_0  (
    .a(\U4/AddrCtrl [0]),
    .b(1'b0),
    .c(\U4/lt2_c0 ),
    .o({\U4/lt2_c1 ,open_n329}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt2_1  (
    .a(\U4/AddrCtrl [1]),
    .b(1'b0),
    .c(\U4/lt2_c1 ),
    .o({\U4/lt2_c2 ,open_n330}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt2_10  (
    .a(\U4/AddrCtrl [10]),
    .b(1'b0),
    .c(\U4/lt2_c10 ),
    .o({\U4/lt2_c11 ,open_n331}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt2_11  (
    .a(\U4/AddrCtrl [11]),
    .b(1'b0),
    .c(\U4/lt2_c11 ),
    .o({\U4/lt2_c12 ,open_n332}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt2_12  (
    .a(\U4/AddrCtrl [12]),
    .b(1'b0),
    .c(\U4/lt2_c12 ),
    .o({\U4/lt2_c13 ,open_n333}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt2_13  (
    .a(\U4/AddrCtrl [13]),
    .b(1'b0),
    .c(\U4/lt2_c13 ),
    .o({\U4/lt2_c14 ,open_n334}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt2_14  (
    .a(\U4/AddrCtrl [14]),
    .b(1'b0),
    .c(\U4/lt2_c14 ),
    .o({\U4/lt2_c15 ,open_n335}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt2_15  (
    .a(\U4/AddrCtrl [15]),
    .b(1'b0),
    .c(\U4/lt2_c15 ),
    .o({\U4/lt2_c16 ,open_n336}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt2_2  (
    .a(\U4/AddrCtrl [2]),
    .b(1'b0),
    .c(\U4/lt2_c2 ),
    .o({\U4/lt2_c3 ,open_n337}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt2_3  (
    .a(\U4/AddrCtrl [3]),
    .b(1'b0),
    .c(\U4/lt2_c3 ),
    .o({\U4/lt2_c4 ,open_n338}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt2_4  (
    .a(\U4/AddrCtrl [4]),
    .b(1'b1),
    .c(\U4/lt2_c4 ),
    .o({\U4/lt2_c5 ,open_n339}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt2_5  (
    .a(\U4/AddrCtrl [5]),
    .b(1'b0),
    .c(\U4/lt2_c5 ),
    .o({\U4/lt2_c6 ,open_n340}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt2_6  (
    .a(\U4/AddrCtrl [6]),
    .b(1'b0),
    .c(\U4/lt2_c6 ),
    .o({\U4/lt2_c7 ,open_n341}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt2_7  (
    .a(\U4/AddrCtrl [7]),
    .b(1'b1),
    .c(\U4/lt2_c7 ),
    .o({\U4/lt2_c8 ,open_n342}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt2_8  (
    .a(\U4/AddrCtrl [8]),
    .b(1'b1),
    .c(\U4/lt2_c8 ),
    .o({\U4/lt2_c9 ,open_n343}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt2_9  (
    .a(\U4/AddrCtrl [9]),
    .b(1'b0),
    .c(\U4/lt2_c9 ),
    .o({\U4/lt2_c10 ,open_n344}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \U4/lt2_cin  (
    .a(1'b0),
    .o({\U4/lt2_c0 ,open_n347}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt2_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\U4/lt2_c16 ),
    .o({open_n348,\U4/n27 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt3_0  (
    .a(1'b0),
    .b(\U4/AddrCtrl [0]),
    .c(\U4/lt3_c0 ),
    .o({\U4/lt3_c1 ,open_n349}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt3_1  (
    .a(1'b0),
    .b(\U4/AddrCtrl [1]),
    .c(\U4/lt3_c1 ),
    .o({\U4/lt3_c2 ,open_n350}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt3_10  (
    .a(1'b0),
    .b(\U4/AddrCtrl [10]),
    .c(\U4/lt3_c10 ),
    .o({\U4/lt3_c11 ,open_n351}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt3_11  (
    .a(1'b0),
    .b(\U4/AddrCtrl [11]),
    .c(\U4/lt3_c11 ),
    .o({\U4/lt3_c12 ,open_n352}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt3_12  (
    .a(1'b0),
    .b(\U4/AddrCtrl [12]),
    .c(\U4/lt3_c12 ),
    .o({\U4/lt3_c13 ,open_n353}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt3_13  (
    .a(1'b0),
    .b(\U4/AddrCtrl [13]),
    .c(\U4/lt3_c13 ),
    .o({\U4/lt3_c14 ,open_n354}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt3_14  (
    .a(1'b0),
    .b(\U4/AddrCtrl [14]),
    .c(\U4/lt3_c14 ),
    .o({\U4/lt3_c15 ,open_n355}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt3_15  (
    .a(1'b0),
    .b(\U4/AddrCtrl [15]),
    .c(\U4/lt3_c15 ),
    .o({\U4/lt3_c16 ,open_n356}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt3_2  (
    .a(1'b0),
    .b(\U4/AddrCtrl [2]),
    .c(\U4/lt3_c2 ),
    .o({\U4/lt3_c3 ,open_n357}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt3_3  (
    .a(1'b0),
    .b(\U4/AddrCtrl [3]),
    .c(\U4/lt3_c3 ),
    .o({\U4/lt3_c4 ,open_n358}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt3_4  (
    .a(1'b1),
    .b(\U4/AddrCtrl [4]),
    .c(\U4/lt3_c4 ),
    .o({\U4/lt3_c5 ,open_n359}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt3_5  (
    .a(1'b0),
    .b(\U4/AddrCtrl [5]),
    .c(\U4/lt3_c5 ),
    .o({\U4/lt3_c6 ,open_n360}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt3_6  (
    .a(1'b0),
    .b(\U4/AddrCtrl [6]),
    .c(\U4/lt3_c6 ),
    .o({\U4/lt3_c7 ,open_n361}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt3_7  (
    .a(1'b1),
    .b(\U4/AddrCtrl [7]),
    .c(\U4/lt3_c7 ),
    .o({\U4/lt3_c8 ,open_n362}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt3_8  (
    .a(1'b1),
    .b(\U4/AddrCtrl [8]),
    .c(\U4/lt3_c8 ),
    .o({\U4/lt3_c9 ,open_n363}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt3_9  (
    .a(1'b0),
    .b(\U4/AddrCtrl [9]),
    .c(\U4/lt3_c9 ),
    .o({\U4/lt3_c10 ,open_n364}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \U4/lt3_cin  (
    .a(1'b1),
    .o({\U4/lt3_c0 ,open_n367}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt3_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\U4/lt3_c16 ),
    .o({open_n368,\U4/n31 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt4_0  (
    .a(\U4/AddrCtrl [0]),
    .b(1'b0),
    .c(\U4/lt4_c0 ),
    .o({\U4/lt4_c1 ,open_n369}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt4_1  (
    .a(\U4/AddrCtrl [1]),
    .b(1'b0),
    .c(\U4/lt4_c1 ),
    .o({\U4/lt4_c2 ,open_n370}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt4_10  (
    .a(\U4/AddrCtrl [10]),
    .b(1'b0),
    .c(\U4/lt4_c10 ),
    .o({\U4/lt4_c11 ,open_n371}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt4_11  (
    .a(\U4/AddrCtrl [11]),
    .b(1'b0),
    .c(\U4/lt4_c11 ),
    .o({\U4/lt4_c12 ,open_n372}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt4_12  (
    .a(\U4/AddrCtrl [12]),
    .b(1'b0),
    .c(\U4/lt4_c12 ),
    .o({\U4/lt4_c13 ,open_n373}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt4_13  (
    .a(\U4/AddrCtrl [13]),
    .b(1'b0),
    .c(\U4/lt4_c13 ),
    .o({\U4/lt4_c14 ,open_n374}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt4_14  (
    .a(\U4/AddrCtrl [14]),
    .b(1'b0),
    .c(\U4/lt4_c14 ),
    .o({\U4/lt4_c15 ,open_n375}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt4_15  (
    .a(\U4/AddrCtrl [15]),
    .b(1'b0),
    .c(\U4/lt4_c15 ),
    .o({\U4/lt4_c16 ,open_n376}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt4_2  (
    .a(\U4/AddrCtrl [2]),
    .b(1'b0),
    .c(\U4/lt4_c2 ),
    .o({\U4/lt4_c3 ,open_n377}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt4_3  (
    .a(\U4/AddrCtrl [3]),
    .b(1'b0),
    .c(\U4/lt4_c3 ),
    .o({\U4/lt4_c4 ,open_n378}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt4_4  (
    .a(\U4/AddrCtrl [4]),
    .b(1'b0),
    .c(\U4/lt4_c4 ),
    .o({\U4/lt4_c5 ,open_n379}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt4_5  (
    .a(\U4/AddrCtrl [5]),
    .b(1'b1),
    .c(\U4/lt4_c5 ),
    .o({\U4/lt4_c6 ,open_n380}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt4_6  (
    .a(\U4/AddrCtrl [6]),
    .b(1'b0),
    .c(\U4/lt4_c6 ),
    .o({\U4/lt4_c7 ,open_n381}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt4_7  (
    .a(\U4/AddrCtrl [7]),
    .b(1'b0),
    .c(\U4/lt4_c7 ),
    .o({\U4/lt4_c8 ,open_n382}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt4_8  (
    .a(\U4/AddrCtrl [8]),
    .b(1'b1),
    .c(\U4/lt4_c8 ),
    .o({\U4/lt4_c9 ,open_n383}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt4_9  (
    .a(\U4/AddrCtrl [9]),
    .b(1'b1),
    .c(\U4/lt4_c9 ),
    .o({\U4/lt4_c10 ,open_n384}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \U4/lt4_cin  (
    .a(1'b0),
    .o({\U4/lt4_c0 ,open_n387}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt4_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\U4/lt4_c16 ),
    .o({open_n388,\U4/n33 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt5_0  (
    .a(1'b0),
    .b(\U4/AddrCtrl [0]),
    .c(\U4/lt5_c0 ),
    .o({\U4/lt5_c1 ,open_n389}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt5_1  (
    .a(1'b0),
    .b(\U4/AddrCtrl [1]),
    .c(\U4/lt5_c1 ),
    .o({\U4/lt5_c2 ,open_n390}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt5_10  (
    .a(1'b0),
    .b(\U4/AddrCtrl [10]),
    .c(\U4/lt5_c10 ),
    .o({\U4/lt5_c11 ,open_n391}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt5_11  (
    .a(1'b0),
    .b(\U4/AddrCtrl [11]),
    .c(\U4/lt5_c11 ),
    .o({\U4/lt5_c12 ,open_n392}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt5_12  (
    .a(1'b0),
    .b(\U4/AddrCtrl [12]),
    .c(\U4/lt5_c12 ),
    .o({\U4/lt5_c13 ,open_n393}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt5_13  (
    .a(1'b0),
    .b(\U4/AddrCtrl [13]),
    .c(\U4/lt5_c13 ),
    .o({\U4/lt5_c14 ,open_n394}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt5_14  (
    .a(1'b0),
    .b(\U4/AddrCtrl [14]),
    .c(\U4/lt5_c14 ),
    .o({\U4/lt5_c15 ,open_n395}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt5_15  (
    .a(1'b0),
    .b(\U4/AddrCtrl [15]),
    .c(\U4/lt5_c15 ),
    .o({\U4/lt5_c16 ,open_n396}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt5_2  (
    .a(1'b0),
    .b(\U4/AddrCtrl [2]),
    .c(\U4/lt5_c2 ),
    .o({\U4/lt5_c3 ,open_n397}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt5_3  (
    .a(1'b0),
    .b(\U4/AddrCtrl [3]),
    .c(\U4/lt5_c3 ),
    .o({\U4/lt5_c4 ,open_n398}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt5_4  (
    .a(1'b0),
    .b(\U4/AddrCtrl [4]),
    .c(\U4/lt5_c4 ),
    .o({\U4/lt5_c5 ,open_n399}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt5_5  (
    .a(1'b1),
    .b(\U4/AddrCtrl [5]),
    .c(\U4/lt5_c5 ),
    .o({\U4/lt5_c6 ,open_n400}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt5_6  (
    .a(1'b0),
    .b(\U4/AddrCtrl [6]),
    .c(\U4/lt5_c6 ),
    .o({\U4/lt5_c7 ,open_n401}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt5_7  (
    .a(1'b0),
    .b(\U4/AddrCtrl [7]),
    .c(\U4/lt5_c7 ),
    .o({\U4/lt5_c8 ,open_n402}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt5_8  (
    .a(1'b1),
    .b(\U4/AddrCtrl [8]),
    .c(\U4/lt5_c8 ),
    .o({\U4/lt5_c9 ,open_n403}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt5_9  (
    .a(1'b1),
    .b(\U4/AddrCtrl [9]),
    .c(\U4/lt5_c9 ),
    .o({\U4/lt5_c10 ,open_n404}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \U4/lt5_cin  (
    .a(1'b1),
    .o({\U4/lt5_c0 ,open_n407}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt5_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\U4/lt5_c16 ),
    .o({open_n408,\U4/n37 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt6_0  (
    .a(\U4/AddrCtrl [0]),
    .b(1'b0),
    .c(\U4/lt6_c0 ),
    .o({\U4/lt6_c1 ,open_n409}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt6_1  (
    .a(\U4/AddrCtrl [1]),
    .b(1'b0),
    .c(\U4/lt6_c1 ),
    .o({\U4/lt6_c2 ,open_n410}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt6_10  (
    .a(\U4/AddrCtrl [10]),
    .b(1'b1),
    .c(\U4/lt6_c10 ),
    .o({\U4/lt6_c11 ,open_n411}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt6_11  (
    .a(\U4/AddrCtrl [11]),
    .b(1'b0),
    .c(\U4/lt6_c11 ),
    .o({\U4/lt6_c12 ,open_n412}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt6_12  (
    .a(\U4/AddrCtrl [12]),
    .b(1'b0),
    .c(\U4/lt6_c12 ),
    .o({\U4/lt6_c13 ,open_n413}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt6_13  (
    .a(\U4/AddrCtrl [13]),
    .b(1'b0),
    .c(\U4/lt6_c13 ),
    .o({\U4/lt6_c14 ,open_n414}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt6_14  (
    .a(\U4/AddrCtrl [14]),
    .b(1'b0),
    .c(\U4/lt6_c14 ),
    .o({\U4/lt6_c15 ,open_n415}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt6_15  (
    .a(\U4/AddrCtrl [15]),
    .b(1'b0),
    .c(\U4/lt6_c15 ),
    .o({\U4/lt6_c16 ,open_n416}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt6_2  (
    .a(\U4/AddrCtrl [2]),
    .b(1'b0),
    .c(\U4/lt6_c2 ),
    .o({\U4/lt6_c3 ,open_n417}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt6_3  (
    .a(\U4/AddrCtrl [3]),
    .b(1'b0),
    .c(\U4/lt6_c3 ),
    .o({\U4/lt6_c4 ,open_n418}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt6_4  (
    .a(\U4/AddrCtrl [4]),
    .b(1'b1),
    .c(\U4/lt6_c4 ),
    .o({\U4/lt6_c5 ,open_n419}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt6_5  (
    .a(\U4/AddrCtrl [5]),
    .b(1'b1),
    .c(\U4/lt6_c5 ),
    .o({\U4/lt6_c6 ,open_n420}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt6_6  (
    .a(\U4/AddrCtrl [6]),
    .b(1'b0),
    .c(\U4/lt6_c6 ),
    .o({\U4/lt6_c7 ,open_n421}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt6_7  (
    .a(\U4/AddrCtrl [7]),
    .b(1'b1),
    .c(\U4/lt6_c7 ),
    .o({\U4/lt6_c8 ,open_n422}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt6_8  (
    .a(\U4/AddrCtrl [8]),
    .b(1'b0),
    .c(\U4/lt6_c8 ),
    .o({\U4/lt6_c9 ,open_n423}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt6_9  (
    .a(\U4/AddrCtrl [9]),
    .b(1'b0),
    .c(\U4/lt6_c9 ),
    .o({\U4/lt6_c10 ,open_n424}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \U4/lt6_cin  (
    .a(1'b0),
    .o({\U4/lt6_c0 ,open_n427}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt6_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\U4/lt6_c16 ),
    .o({open_n428,\U4/n39 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt7_0  (
    .a(1'b0),
    .b(\U4/AddrCtrl [0]),
    .c(\U4/lt7_c0 ),
    .o({\U4/lt7_c1 ,open_n429}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt7_1  (
    .a(1'b0),
    .b(\U4/AddrCtrl [1]),
    .c(\U4/lt7_c1 ),
    .o({\U4/lt7_c2 ,open_n430}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt7_10  (
    .a(1'b1),
    .b(\U4/AddrCtrl [10]),
    .c(\U4/lt7_c10 ),
    .o({\U4/lt7_c11 ,open_n431}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt7_11  (
    .a(1'b0),
    .b(\U4/AddrCtrl [11]),
    .c(\U4/lt7_c11 ),
    .o({\U4/lt7_c12 ,open_n432}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt7_12  (
    .a(1'b0),
    .b(\U4/AddrCtrl [12]),
    .c(\U4/lt7_c12 ),
    .o({\U4/lt7_c13 ,open_n433}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt7_13  (
    .a(1'b0),
    .b(\U4/AddrCtrl [13]),
    .c(\U4/lt7_c13 ),
    .o({\U4/lt7_c14 ,open_n434}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt7_14  (
    .a(1'b0),
    .b(\U4/AddrCtrl [14]),
    .c(\U4/lt7_c14 ),
    .o({\U4/lt7_c15 ,open_n435}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt7_15  (
    .a(1'b0),
    .b(\U4/AddrCtrl [15]),
    .c(\U4/lt7_c15 ),
    .o({\U4/lt7_c16 ,open_n436}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt7_2  (
    .a(1'b0),
    .b(\U4/AddrCtrl [2]),
    .c(\U4/lt7_c2 ),
    .o({\U4/lt7_c3 ,open_n437}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt7_3  (
    .a(1'b0),
    .b(\U4/AddrCtrl [3]),
    .c(\U4/lt7_c3 ),
    .o({\U4/lt7_c4 ,open_n438}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt7_4  (
    .a(1'b1),
    .b(\U4/AddrCtrl [4]),
    .c(\U4/lt7_c4 ),
    .o({\U4/lt7_c5 ,open_n439}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt7_5  (
    .a(1'b1),
    .b(\U4/AddrCtrl [5]),
    .c(\U4/lt7_c5 ),
    .o({\U4/lt7_c6 ,open_n440}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt7_6  (
    .a(1'b0),
    .b(\U4/AddrCtrl [6]),
    .c(\U4/lt7_c6 ),
    .o({\U4/lt7_c7 ,open_n441}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt7_7  (
    .a(1'b1),
    .b(\U4/AddrCtrl [7]),
    .c(\U4/lt7_c7 ),
    .o({\U4/lt7_c8 ,open_n442}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt7_8  (
    .a(1'b0),
    .b(\U4/AddrCtrl [8]),
    .c(\U4/lt7_c8 ),
    .o({\U4/lt7_c9 ,open_n443}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt7_9  (
    .a(1'b0),
    .b(\U4/AddrCtrl [9]),
    .c(\U4/lt7_c9 ),
    .o({\U4/lt7_c10 ,open_n444}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \U4/lt7_cin  (
    .a(1'b1),
    .o({\U4/lt7_c0 ,open_n447}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \U4/lt7_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\U4/lt7_c16 ),
    .o({open_n448,\U4/n43 }));
  reg_ar_as_w1 \U4/reg0_b0  (
    .clk(i8080_WR_pad),
    .d(i8080_D_pad[0]),
    .en(\U4/mux1_b0_sel_is_3_o ),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U4/LCD_Pix_Reg [0]));  // source/LCD8080Ctrl.v(70)
  EF2_PHY_SPAD #(
    //.CLKSRC("CLK"),
    //.LOCATION("P9"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DO_DFFMODE("FF"),
    .DO_REGSET("SET"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .OUTCEMUX("CE"),
    .OUTCLKMUX("CLK"),
    .OUTRSTMUX("INV"),
    .SRMODE("ASYNC"),
    .TSMUX("INV"))
    \U4/reg1_b0_DO  (
    .ce(\U4/mux2_b0_sel_is_3_o ),
    .clk(i8080_WR_pad),
    .do({open_n449,i8080_D_pad[0]}),
    .rst(nRST_pad),
    .ts(1'b1),
    .opad(LCDBK));  // source/LCD8080Ctrl.v(70)
  reg_ar_as_w1 \U4/reg2_b0  (
    .clk(CLK_100M),
    .d(\U4/n21 [0]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U4/AddrCtrl [0]));  // source/LCD8080Ctrl.v(104)
  reg_ar_as_w1 \U4/reg2_b1  (
    .clk(CLK_100M),
    .d(\U4/n21 [1]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U4/AddrCtrl [1]));  // source/LCD8080Ctrl.v(104)
  reg_ar_as_w1 \U4/reg2_b10  (
    .clk(CLK_100M),
    .d(\U4/n21 [10]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U4/AddrCtrl [10]));  // source/LCD8080Ctrl.v(104)
  reg_ar_as_w1 \U4/reg2_b11  (
    .clk(CLK_100M),
    .d(\U4/n21 [11]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U4/AddrCtrl [11]));  // source/LCD8080Ctrl.v(104)
  reg_ar_as_w1 \U4/reg2_b12  (
    .clk(CLK_100M),
    .d(\U4/n21 [12]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U4/AddrCtrl [12]));  // source/LCD8080Ctrl.v(104)
  reg_ar_as_w1 \U4/reg2_b13  (
    .clk(CLK_100M),
    .d(\U4/n21 [13]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U4/AddrCtrl [13]));  // source/LCD8080Ctrl.v(104)
  reg_ar_as_w1 \U4/reg2_b14  (
    .clk(CLK_100M),
    .d(\U4/n21 [14]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U4/AddrCtrl [14]));  // source/LCD8080Ctrl.v(104)
  reg_ar_as_w1 \U4/reg2_b15  (
    .clk(CLK_100M),
    .d(\U4/n21 [15]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U4/AddrCtrl [15]));  // source/LCD8080Ctrl.v(104)
  reg_ar_as_w1 \U4/reg2_b2  (
    .clk(CLK_100M),
    .d(\U4/n21 [2]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U4/AddrCtrl [2]));  // source/LCD8080Ctrl.v(104)
  reg_ar_as_w1 \U4/reg2_b3  (
    .clk(CLK_100M),
    .d(\U4/n21 [3]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U4/AddrCtrl [3]));  // source/LCD8080Ctrl.v(104)
  reg_ar_as_w1 \U4/reg2_b4  (
    .clk(CLK_100M),
    .d(\U4/n21 [4]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U4/AddrCtrl [4]));  // source/LCD8080Ctrl.v(104)
  reg_ar_as_w1 \U4/reg2_b5  (
    .clk(CLK_100M),
    .d(\U4/n21 [5]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U4/AddrCtrl [5]));  // source/LCD8080Ctrl.v(104)
  reg_ar_as_w1 \U4/reg2_b6  (
    .clk(CLK_100M),
    .d(\U4/n21 [6]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U4/AddrCtrl [6]));  // source/LCD8080Ctrl.v(104)
  reg_ar_as_w1 \U4/reg2_b7  (
    .clk(CLK_100M),
    .d(\U4/n21 [7]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U4/AddrCtrl [7]));  // source/LCD8080Ctrl.v(104)
  reg_ar_as_w1 \U4/reg2_b8  (
    .clk(CLK_100M),
    .d(\U4/n21 [8]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U4/AddrCtrl [8]));  // source/LCD8080Ctrl.v(104)
  reg_ar_as_w1 \U4/reg2_b9  (
    .clk(CLK_100M),
    .d(\U4/n21 [9]),
    .en(1'b1),
    .reset(~nRST_pad),
    .set(1'b0),
    .q(\U4/AddrCtrl [9]));  // source/LCD8080Ctrl.v(104)
  EF2_PHY_SPAD #(
    //.CLKSRC("CLK"),
    //.LOCATION("P20"),
    //.PULLMODE("PULLUP"),
    .INCEMUX("CE"),
    .INCLKMUX("CLK"),
    .INRSTMUX("INV"),
    .IN_DFFMODE("FF"),
    .IN_REGSET("SET"),
    .IOTYPE("LVCMOS18"),
    .MODE("IN"),
    .SRMODE("ASYNC"),
    .TSMUX("TS"))
    \U4/reg3_b3_IN  (
    .ce(\U4/mux0_b3_sel_is_3_o ),
    .clk(i8080_WR_pad),
    .ipad(i8080_D[3]),
    .rst(nRST_pad),
    .ts(1'b1),
    .di(i8080_D_pad[3]),
    .diq({open_n457,\U4/LCD_Ctrl_Reg [3]}));  // source/LCD8080Ctrl.v(70)
  EF2_PHY_SPAD #(
    //.CLKSRC("CLK"),
    //.LOCATION("P19"),
    //.PULLMODE("PULLUP"),
    .INCEMUX("CE"),
    .INCLKMUX("CLK"),
    .INRSTMUX("INV"),
    .IN_DFFMODE("FF"),
    .IN_REGSET("RESET"),
    .IOTYPE("LVCMOS18"),
    .MODE("IN"),
    .SRMODE("ASYNC"),
    .TSMUX("TS"))
    \U4/reg3_b4_IN  (
    .ce(\U4/mux0_b3_sel_is_3_o ),
    .clk(i8080_WR_pad),
    .ipad(i8080_D[4]),
    .rst(nRST_pad),
    .ts(1'b1),
    .di(i8080_D_pad[4]),
    .diq({open_n462,\U4/LCD_Ctrl_Reg [4]}));  // source/LCD8080Ctrl.v(70)
  EF2_PHY_SPAD #(
    //.LOCATION("P24"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS18"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u100 (
    .ipad(i8080_D[1]),
    .ts(1'b1),
    .di(i8080_D_pad[1]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(12)
  EF2_PHY_SPAD #(
    //.LOCATION("P25"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS18"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u101 (
    .ipad(i8080_D[0]),
    .ts(1'b1),
    .di(i8080_D_pad[0]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(12)
  EF2_PHY_SPAD #(
    //.LOCATION("P13"),
    //.PULLMODE("PULLUP"),
    //.SLEWRATE("MED"),
    .DRIVE("12"),
    .IOTYPE("LVCMOS18"),
    .MODE("BI"),
    .TO_DFFMODE("NONE"),
    .TSMUX("INV"))
    _al_u102 (
    .do({open_n485,\U4/FrameSync }),
    .ts(\U4/LCD_Ctrl_Reg [4]),
    .di(i8080_RS_pad),
    .bpad(i8080_RS));  // source/LCD8080Ctrl.v(73)
  EF2_PHY_SPAD #(
    //.LOCATION("P14"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS18"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u103 (
    .ipad(i8080_WR),
    .ts(1'b1),
    .di(i8080_WR_pad));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(10)
  EF2_PHY_SPAD #(
    //.LOCATION("P12"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u104 (
    .ipad(nRST),
    .ts(1'b1),
    .di(nRST_pad));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(4)
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u107 (
    .a(FIFO_EMPTY),
    .b(FIFO_DO[3]),
    .o(LCD_B_pad[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u108 (
    .a(FIFO_EMPTY),
    .b(FIFO_DO[2]),
    .o(LCD_B_pad[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u109 (
    .a(FIFO_EMPTY),
    .b(FIFO_DO[1]),
    .o(LCD_B_pad[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u110 (
    .a(FIFO_EMPTY),
    .b(FIFO_DO[0]),
    .o(LCD_B_pad[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u111 (
    .a(FIFO_EMPTY),
    .b(FIFO_DO[10]),
    .o(LCD_G_pad[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u112 (
    .a(FIFO_EMPTY),
    .b(FIFO_DO[9]),
    .o(LCD_G_pad[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u113 (
    .a(FIFO_EMPTY),
    .b(FIFO_DO[8]),
    .o(LCD_G_pad[5]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u114 (
    .a(FIFO_DO[11]),
    .b(FIFO_EMPTY),
    .o(LCD_R_pad[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u115 (
    .a(FIFO_EMPTY),
    .b(FIFO_DO[7]),
    .o(LCD_G_pad[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u116 (
    .a(FIFO_EMPTY),
    .b(FIFO_DO[6]),
    .o(LCD_G_pad[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u117 (
    .a(FIFO_EMPTY),
    .b(FIFO_DO[5]),
    .o(LCD_G_pad[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u118 (
    .a(FIFO_EMPTY),
    .b(FIFO_DO[4]),
    .o(LCD_B_pad[7]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u119 (
    .a(FIFO_EMPTY),
    .b(FIFO_DO[15]),
    .o(LCD_R_pad[7]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u120 (
    .a(FIFO_EMPTY),
    .b(FIFO_DO[14]),
    .o(LCD_R_pad[6]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u121 (
    .a(FIFO_EMPTY),
    .b(FIFO_DO[13]),
    .o(LCD_R_pad[5]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u122 (
    .a(FIFO_EMPTY),
    .b(FIFO_DO[12]),
    .o(LCD_R_pad[4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u123 (
    .a(CLK_100M),
    .b(i8080_WR_pad),
    .c(\U4/LCD_Ctrl_Reg [4]),
    .o(FIFO_CLK_W));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u124 (
    .a(\D1/n14 ),
    .b(\D1/n15 ),
    .o(LCD_HYNC_pad));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u125 (
    .a(LCD_HYNC_pad),
    .b(LCD_SYNC_pad),
    .o(_al_u125_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u126 (
    .a(\U4/n18 [9]),
    .b(\U4/AddrCtrl [9]),
    .c(\U4/n17 ),
    .d(_al_u125_o),
    .o(\U4/n21 [9]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u127 (
    .a(\U4/n18 [8]),
    .b(\U4/AddrCtrl [8]),
    .c(\U4/n17 ),
    .d(_al_u125_o),
    .o(\U4/n21 [8]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u128 (
    .a(\U4/n18 [7]),
    .b(\U4/AddrCtrl [7]),
    .c(\U4/n17 ),
    .d(_al_u125_o),
    .o(\U4/n21 [7]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u129 (
    .a(\U4/n18 [6]),
    .b(\U4/AddrCtrl [6]),
    .c(\U4/n17 ),
    .d(_al_u125_o),
    .o(\U4/n21 [6]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u130 (
    .a(\U4/n18 [5]),
    .b(\U4/AddrCtrl [5]),
    .c(\U4/n17 ),
    .d(_al_u125_o),
    .o(\U4/n21 [5]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u131 (
    .a(\U4/n18 [4]),
    .b(\U4/AddrCtrl [4]),
    .c(\U4/n17 ),
    .d(_al_u125_o),
    .o(\U4/n21 [4]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u132 (
    .a(\U4/n18 [3]),
    .b(\U4/AddrCtrl [3]),
    .c(\U4/n17 ),
    .d(_al_u125_o),
    .o(\U4/n21 [3]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u133 (
    .a(\U4/n18 [2]),
    .b(\U4/AddrCtrl [2]),
    .c(\U4/n17 ),
    .d(_al_u125_o),
    .o(\U4/n21 [2]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u134 (
    .a(\U4/n18 [1]),
    .b(\U4/AddrCtrl [1]),
    .c(\U4/n17 ),
    .d(_al_u125_o),
    .o(\U4/n21 [1]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u135 (
    .a(\U4/n18 [15]),
    .b(\U4/AddrCtrl [15]),
    .c(\U4/n17 ),
    .d(_al_u125_o),
    .o(\U4/n21 [15]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u136 (
    .a(\U4/n18 [14]),
    .b(\U4/AddrCtrl [14]),
    .c(\U4/n17 ),
    .d(_al_u125_o),
    .o(\U4/n21 [14]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u137 (
    .a(\U4/n18 [13]),
    .b(\U4/AddrCtrl [13]),
    .c(\U4/n17 ),
    .d(_al_u125_o),
    .o(\U4/n21 [13]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u138 (
    .a(\U4/n18 [12]),
    .b(\U4/AddrCtrl [12]),
    .c(\U4/n17 ),
    .d(_al_u125_o),
    .o(\U4/n21 [12]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u139 (
    .a(\U4/n18 [11]),
    .b(\U4/AddrCtrl [11]),
    .c(\U4/n17 ),
    .d(_al_u125_o),
    .o(\U4/n21 [11]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u140 (
    .a(\U4/n18 [10]),
    .b(\U4/AddrCtrl [10]),
    .c(\U4/n17 ),
    .d(_al_u125_o),
    .o(\U4/n21 [10]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u141 (
    .a(\U4/n18 [0]),
    .b(\U4/AddrCtrl [0]),
    .c(\U4/n17 ),
    .d(_al_u125_o),
    .o(\U4/n21 [0]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u142 (
    .a(\D1/n17 ),
    .b(\D1/n18 ),
    .c(\D1/n20 ),
    .d(\D1/n22 ),
    .o(LCD_DEN_pad));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u143 (
    .a(LCD_HYNC_pad),
    .b(\U4/LCD_Ctrl_Reg [3]),
    .c(LCD_SYNC_pad),
    .o(\U4/FrameSync ));
  AL_MAP_LUT4 #(
    .EQN("~(~(B*A)*~(C)*~(D)+~(B*A)*C*~(D)+~(~(B*A))*C*D+~(B*A)*C*D)"),
    .INIT(16'h0f88))
    _al_u144 (
    .a(_al_u125_o),
    .b(\U4/n23 ),
    .c(i8080_CS_pad),
    .d(\U4/LCD_Ctrl_Reg [4]),
    .o(FIFO_WE));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*~A)"),
    .INIT(32'h40000000))
    _al_u145 (
    .a(FIFO_EMPTY),
    .b(\D1/n22 ),
    .c(\D1/n24 ),
    .d(\D1/n26 ),
    .e(\D1/n20 ),
    .o(FIFO_RE));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~C*~B*~A)"),
    .INIT(32'h01000000))
    _al_u146 (
    .a(i8080_CS_pad),
    .b(i8080_D_pad[7]),
    .c(i8080_D_pad[6]),
    .d(i8080_RS_pad),
    .e(i8080_D_pad[5]),
    .o(\U4/mux0_b3_sel_is_3_o ));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*~B*~A)"),
    .INIT(32'h10000000))
    _al_u147 (
    .a(i8080_CS_pad),
    .b(i8080_D_pad[7]),
    .c(i8080_RS_pad),
    .d(i8080_D_pad[6]),
    .e(i8080_D_pad[5]),
    .o(\U4/mux2_b0_sel_is_3_o ));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~C*~B*~A)"),
    .INIT(32'h01000000))
    _al_u148 (
    .a(i8080_CS_pad),
    .b(i8080_D_pad[7]),
    .c(i8080_D_pad[5]),
    .d(i8080_D_pad[6]),
    .e(i8080_RS_pad),
    .o(\U4/mux1_b0_sel_is_3_o ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u149 (
    .a(\D1/LineCount [0]),
    .b(\D1/LineCount [1]),
    .c(\D1/LineCount [10]),
    .d(\D1/LineCount [11]),
    .o(_al_u149_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*~A)"),
    .INIT(32'h00010000))
    _al_u150 (
    .a(\D1/LineCount [12]),
    .b(\D1/LineCount [13]),
    .c(\D1/LineCount [14]),
    .d(\D1/LineCount [15]),
    .e(_al_u149_o),
    .o(_al_u150_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*~A)"),
    .INIT(16'h1000))
    _al_u151 (
    .a(\D1/LineCount [3]),
    .b(\D1/LineCount [4]),
    .c(\D1/LineCount [2]),
    .d(\D1/LineCount [5]),
    .o(_al_u151_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~C*~B*~A)"),
    .INIT(32'h01000000))
    _al_u152 (
    .a(\D1/LineCount [6]),
    .b(\D1/LineCount [7]),
    .c(\D1/LineCount [9]),
    .d(\D1/LineCount [8]),
    .e(_al_u151_o),
    .o(_al_u152_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u153 (
    .a(_al_u150_o),
    .b(_al_u152_o),
    .o(_al_u153_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~B*~A))"),
    .INIT(16'h00fe))
    _al_u154 (
    .a(\U4/LCD_Pix_Reg [0]),
    .b(\U4/LCD_Ctrl_Reg [3]),
    .c(\D1/FrameFlag ),
    .d(_al_u153_o),
    .o(\D1/n13 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*~A)"),
    .INIT(16'h1000))
    _al_u155 (
    .a(\U1/Count [25]),
    .b(\U1/Count [26]),
    .c(\U1/Count [23]),
    .d(\U1/Count [24]),
    .o(_al_u155_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*~A)"),
    .INIT(32'h00010000))
    _al_u156 (
    .a(\U1/Count [27]),
    .b(\U1/Count [28]),
    .c(\U1/Count [29]),
    .d(\U1/Count [3]),
    .e(_al_u155_o),
    .o(_al_u156_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u157 (
    .a(\U1/Count [30]),
    .b(\U1/Count [31]),
    .c(\U1/Count [4]),
    .d(\U1/Count [5]),
    .o(_al_u157_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*~B*~A)"),
    .INIT(32'h10000000))
    _al_u158 (
    .a(\U1/Count [7]),
    .b(\U1/Count [8]),
    .c(_al_u157_o),
    .d(\U1/Count [6]),
    .e(\U1/Count [9]),
    .o(_al_u158_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u159 (
    .a(\U1/Count [0]),
    .b(\U1/Count [1]),
    .c(\U1/Count [10]),
    .d(\U1/Count [11]),
    .o(_al_u159_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~C*~B*~A)"),
    .INIT(32'h01000000))
    _al_u160 (
    .a(\U1/Count [12]),
    .b(\U1/Count [13]),
    .c(\U1/Count [14]),
    .d(_al_u159_o),
    .e(\U1/Count [15]),
    .o(_al_u160_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u161 (
    .a(\U1/Count [19]),
    .b(\U1/Count [17]),
    .c(\U1/Count [18]),
    .d(\U1/Count [16]),
    .o(_al_u161_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*~A)"),
    .INIT(32'h40000000))
    _al_u162 (
    .a(\U1/Count [2]),
    .b(_al_u161_o),
    .c(\U1/Count [20]),
    .d(\U1/Count [21]),
    .e(\U1/Count [22]),
    .o(_al_u162_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u163 (
    .a(_al_u156_o),
    .b(_al_u158_o),
    .c(_al_u160_o),
    .d(_al_u162_o),
    .o(\U1/n1 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u164 (
    .a(\U2/Count [23]),
    .b(\U2/Count [25]),
    .c(\U2/Count [26]),
    .d(\U2/Count [24]),
    .o(_al_u164_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*~A)"),
    .INIT(32'h00010000))
    _al_u165 (
    .a(\U2/Count [27]),
    .b(\U2/Count [28]),
    .c(\U2/Count [29]),
    .d(\U2/Count [3]),
    .e(_al_u164_o),
    .o(_al_u165_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u166 (
    .a(\U2/Count [30]),
    .b(\U2/Count [31]),
    .c(\U2/Count [4]),
    .d(\U2/Count [5]),
    .o(_al_u166_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~C*~B*~A)"),
    .INIT(32'h01000000))
    _al_u167 (
    .a(\U2/Count [7]),
    .b(\U2/Count [8]),
    .c(\U2/Count [9]),
    .d(\U2/Count [6]),
    .e(_al_u166_o),
    .o(_al_u167_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u168 (
    .a(\U2/Count [0]),
    .b(\U2/Count [1]),
    .c(\U2/Count [10]),
    .d(\U2/Count [11]),
    .o(_al_u168_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*~A)"),
    .INIT(32'h40000000))
    _al_u169 (
    .a(\U2/Count [15]),
    .b(\U2/Count [12]),
    .c(\U2/Count [13]),
    .d(\U2/Count [14]),
    .e(_al_u168_o),
    .o(_al_u169_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u170 (
    .a(\U2/Count [17]),
    .b(\U2/Count [16]),
    .c(\U2/Count [18]),
    .d(\U2/Count [19]),
    .o(_al_u170_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*~A)"),
    .INIT(32'h40000000))
    _al_u171 (
    .a(\U2/Count [2]),
    .b(_al_u170_o),
    .c(\U2/Count [20]),
    .d(\U2/Count [21]),
    .e(\U2/Count [22]),
    .o(_al_u171_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u172 (
    .a(_al_u165_o),
    .b(_al_u167_o),
    .c(_al_u169_o),
    .d(_al_u171_o),
    .o(\U2/n1 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u173 (
    .a(\D1/PixelCount [0]),
    .b(\D1/PixelCount [1]),
    .c(\D1/PixelCount [10]),
    .d(\D1/PixelCount [11]),
    .o(_al_u173_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*~A)"),
    .INIT(32'h00010000))
    _al_u174 (
    .a(\D1/PixelCount [12]),
    .b(\D1/PixelCount [13]),
    .c(\D1/PixelCount [14]),
    .d(\D1/PixelCount [15]),
    .e(_al_u173_o),
    .o(_al_u174_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u175 (
    .a(\D1/PixelCount [2]),
    .b(\D1/PixelCount [3]),
    .c(\D1/PixelCount [5]),
    .d(\D1/PixelCount [4]),
    .o(_al_u175_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*~A)"),
    .INIT(32'h40000000))
    _al_u176 (
    .a(\D1/PixelCount [8]),
    .b(\D1/PixelCount [6]),
    .c(\D1/PixelCount [7]),
    .d(_al_u175_o),
    .e(\D1/PixelCount [9]),
    .o(_al_u176_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u177 (
    .a(_al_u174_o),
    .b(_al_u176_o),
    .o(_al_u177_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u178 (
    .a(\D1/n2 [9]),
    .b(\D1/LineCount [9]),
    .c(_al_u177_o),
    .o(\D1/n9 [9]));
  AL_MAP_LUT4 #(
    .EQN("((B*~A)*~(C)*~(D)+(B*~A)*C*~(D)+~((B*~A))*C*D+(B*~A)*C*D)"),
    .INIT(16'hf044))
    _al_u179 (
    .a(_al_u153_o),
    .b(\D1/LineCount [8]),
    .c(\D1/n2 [8]),
    .d(_al_u177_o),
    .o(\D1/n9 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u180 (
    .a(\D1/n2 [7]),
    .b(\D1/LineCount [7]),
    .c(_al_u177_o),
    .o(\D1/n9 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u181 (
    .a(\D1/n2 [6]),
    .b(\D1/LineCount [6]),
    .c(_al_u177_o),
    .o(\D1/n9 [6]));
  AL_MAP_LUT4 #(
    .EQN("((B*~A)*~(C)*~(D)+(B*~A)*C*~(D)+~((B*~A))*C*D+(B*~A)*C*D)"),
    .INIT(16'hf044))
    _al_u182 (
    .a(_al_u153_o),
    .b(\D1/LineCount [5]),
    .c(\D1/n2 [5]),
    .d(_al_u177_o),
    .o(\D1/n9 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u183 (
    .a(\D1/n2 [4]),
    .b(\D1/LineCount [4]),
    .c(_al_u177_o),
    .o(\D1/n9 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u184 (
    .a(\D1/n2 [3]),
    .b(\D1/LineCount [3]),
    .c(_al_u177_o),
    .o(\D1/n9 [3]));
  AL_MAP_LUT4 #(
    .EQN("((B*~A)*~(C)*~(D)+(B*~A)*C*~(D)+~((B*~A))*C*D+(B*~A)*C*D)"),
    .INIT(16'hf044))
    _al_u185 (
    .a(_al_u153_o),
    .b(\D1/LineCount [2]),
    .c(\D1/n2 [2]),
    .d(_al_u177_o),
    .o(\D1/n9 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u186 (
    .a(\D1/n2 [15]),
    .b(\D1/LineCount [15]),
    .c(_al_u177_o),
    .o(\D1/n9 [15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u187 (
    .a(\D1/n2 [14]),
    .b(\D1/LineCount [14]),
    .c(_al_u177_o),
    .o(\D1/n9 [14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u188 (
    .a(\D1/n2 [13]),
    .b(\D1/LineCount [13]),
    .c(_al_u177_o),
    .o(\D1/n9 [13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u189 (
    .a(\D1/n2 [12]),
    .b(\D1/LineCount [12]),
    .c(_al_u177_o),
    .o(\D1/n9 [12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u190 (
    .a(\D1/n2 [11]),
    .b(\D1/LineCount [11]),
    .c(_al_u177_o),
    .o(\D1/n9 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u191 (
    .a(\D1/n2 [10]),
    .b(\D1/LineCount [10]),
    .c(_al_u177_o),
    .o(\D1/n9 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u192 (
    .a(\D1/n2 [1]),
    .b(\D1/LineCount [1]),
    .c(_al_u177_o),
    .o(\D1/n9 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u193 (
    .a(\D1/n2 [0]),
    .b(\D1/LineCount [0]),
    .c(_al_u177_o),
    .o(\D1/n9 [0]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u194 (
    .a(\U1/n1 ),
    .b(\U1/n3 [9]),
    .o(\U1/n5 [9]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u195 (
    .a(\U1/n1 ),
    .b(\U1/n3 [8]),
    .o(\U1/n5 [8]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u196 (
    .a(\U1/n1 ),
    .b(\U1/n3 [7]),
    .o(\U1/n5 [7]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u197 (
    .a(\U1/n1 ),
    .b(\U1/n3 [6]),
    .o(\U1/n5 [6]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u198 (
    .a(\U1/n1 ),
    .b(\U1/n3 [5]),
    .o(\U1/n5 [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u199 (
    .a(\U1/n1 ),
    .b(\U1/n3 [4]),
    .o(\U1/n5 [4]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u200 (
    .a(\U1/n1 ),
    .b(\U1/n3 [31]),
    .o(\U1/n5 [31]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u201 (
    .a(\U1/n1 ),
    .b(\U1/n3 [30]),
    .o(\U1/n5 [30]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u202 (
    .a(\U1/n1 ),
    .b(\U1/n3 [3]),
    .o(\U1/n5 [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u203 (
    .a(\U1/n1 ),
    .b(\U1/n3 [29]),
    .o(\U1/n5 [29]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u204 (
    .a(\U1/n1 ),
    .b(\U1/n3 [28]),
    .o(\U1/n5 [28]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u205 (
    .a(\U1/n1 ),
    .b(\U1/n3 [27]),
    .o(\U1/n5 [27]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u206 (
    .a(\U1/n1 ),
    .b(\U1/n3 [26]),
    .o(\U1/n5 [26]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u207 (
    .a(\U1/n1 ),
    .b(\U1/n3 [25]),
    .o(\U1/n5 [25]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u208 (
    .a(\U1/n1 ),
    .b(\U1/n3 [24]),
    .o(\U1/n5 [24]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u209 (
    .a(\U1/n1 ),
    .b(\U1/n3 [23]),
    .o(\U1/n5 [23]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u210 (
    .a(\U1/n1 ),
    .b(\U1/n3 [22]),
    .o(\U1/n5 [22]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u211 (
    .a(\U1/n1 ),
    .b(\U1/n3 [21]),
    .o(\U1/n5 [21]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u212 (
    .a(\U1/n1 ),
    .b(\U1/n3 [20]),
    .o(\U1/n5 [20]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u213 (
    .a(\U1/n1 ),
    .b(\U1/n3 [2]),
    .o(\U1/n5 [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u214 (
    .a(\U1/n1 ),
    .b(\U1/n3 [19]),
    .o(\U1/n5 [19]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u215 (
    .a(\U1/n1 ),
    .b(\U1/n3 [18]),
    .o(\U1/n5 [18]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u216 (
    .a(\U1/n1 ),
    .b(\U1/n3 [17]),
    .o(\U1/n5 [17]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u217 (
    .a(\U1/n1 ),
    .b(\U1/n3 [16]),
    .o(\U1/n5 [16]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u218 (
    .a(\U1/n1 ),
    .b(\U1/n3 [15]),
    .o(\U1/n5 [15]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u219 (
    .a(\U1/n1 ),
    .b(\U1/n3 [14]),
    .o(\U1/n5 [14]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u220 (
    .a(\U1/n1 ),
    .b(\U1/n3 [13]),
    .o(\U1/n5 [13]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u221 (
    .a(\U1/n1 ),
    .b(\U1/n3 [12]),
    .o(\U1/n5 [12]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u222 (
    .a(\U1/n1 ),
    .b(\U1/n3 [11]),
    .o(\U1/n5 [11]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u223 (
    .a(\U1/n1 ),
    .b(\U1/n3 [10]),
    .o(\U1/n5 [10]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u224 (
    .a(\U1/n1 ),
    .b(\U1/n3 [1]),
    .o(\U1/n5 [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u225 (
    .a(\U1/n1 ),
    .b(\U1/n3 [0]),
    .o(\U1/n5 [0]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u226 (
    .a(\U2/n1 ),
    .b(\U2/n3 [9]),
    .o(\U2/n5 [9]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u227 (
    .a(\U2/n1 ),
    .b(\U2/n3 [8]),
    .o(\U2/n5 [8]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u228 (
    .a(\U2/n1 ),
    .b(\U2/n3 [7]),
    .o(\U2/n5 [7]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u229 (
    .a(\U2/n1 ),
    .b(\U2/n3 [6]),
    .o(\U2/n5 [6]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u230 (
    .a(\U2/n1 ),
    .b(\U2/n3 [5]),
    .o(\U2/n5 [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u231 (
    .a(\U2/n1 ),
    .b(\U2/n3 [4]),
    .o(\U2/n5 [4]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u232 (
    .a(\U2/n1 ),
    .b(\U2/n3 [31]),
    .o(\U2/n5 [31]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u233 (
    .a(\U2/n1 ),
    .b(\U2/n3 [30]),
    .o(\U2/n5 [30]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u234 (
    .a(\U2/n1 ),
    .b(\U2/n3 [3]),
    .o(\U2/n5 [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u235 (
    .a(\U2/n1 ),
    .b(\U2/n3 [29]),
    .o(\U2/n5 [29]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u236 (
    .a(\U2/n1 ),
    .b(\U2/n3 [28]),
    .o(\U2/n5 [28]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u237 (
    .a(\U2/n1 ),
    .b(\U2/n3 [27]),
    .o(\U2/n5 [27]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u238 (
    .a(\U2/n1 ),
    .b(\U2/n3 [26]),
    .o(\U2/n5 [26]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u239 (
    .a(\U2/n1 ),
    .b(\U2/n3 [25]),
    .o(\U2/n5 [25]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u240 (
    .a(\U2/n1 ),
    .b(\U2/n3 [24]),
    .o(\U2/n5 [24]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u241 (
    .a(\U2/n1 ),
    .b(\U2/n3 [23]),
    .o(\U2/n5 [23]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u242 (
    .a(\U2/n1 ),
    .b(\U2/n3 [22]),
    .o(\U2/n5 [22]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u243 (
    .a(\U2/n1 ),
    .b(\U2/n3 [21]),
    .o(\U2/n5 [21]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u244 (
    .a(\U2/n1 ),
    .b(\U2/n3 [20]),
    .o(\U2/n5 [20]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u245 (
    .a(\U2/n1 ),
    .b(\U2/n3 [2]),
    .o(\U2/n5 [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u246 (
    .a(\U2/n1 ),
    .b(\U2/n3 [19]),
    .o(\U2/n5 [19]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u247 (
    .a(\U2/n1 ),
    .b(\U2/n3 [18]),
    .o(\U2/n5 [18]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u248 (
    .a(\U2/n1 ),
    .b(\U2/n3 [17]),
    .o(\U2/n5 [17]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u249 (
    .a(\U2/n1 ),
    .b(\U2/n3 [16]),
    .o(\U2/n5 [16]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u250 (
    .a(\U2/n1 ),
    .b(\U2/n3 [15]),
    .o(\U2/n5 [15]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u251 (
    .a(\U2/n1 ),
    .b(\U2/n3 [14]),
    .o(\U2/n5 [14]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u252 (
    .a(\U2/n1 ),
    .b(\U2/n3 [13]),
    .o(\U2/n5 [13]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u253 (
    .a(\U2/n1 ),
    .b(\U2/n3 [12]),
    .o(\U2/n5 [12]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u254 (
    .a(\U2/n1 ),
    .b(\U2/n3 [11]),
    .o(\U2/n5 [11]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u255 (
    .a(\U2/n1 ),
    .b(\U2/n3 [10]),
    .o(\U2/n5 [10]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u256 (
    .a(\U2/n1 ),
    .b(\U2/n3 [1]),
    .o(\U2/n5 [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u257 (
    .a(\U2/n1 ),
    .b(\U2/n3 [0]),
    .o(\U2/n5 [0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u258 (
    .a(_al_u153_o),
    .b(_al_u177_o),
    .o(\D1/mux3_b0_sel_is_0_o ));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u259 (
    .a(\D1/n4 [9]),
    .b(\D1/PixelCount [9]),
    .c(\D1/FrameFlag ),
    .d(\D1/mux3_b0_sel_is_0_o ),
    .o(\D1/n8 [9]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u260 (
    .a(\D1/n4 [8]),
    .b(\D1/PixelCount [8]),
    .c(\D1/FrameFlag ),
    .d(\D1/mux3_b0_sel_is_0_o ),
    .o(\D1/n8 [8]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u261 (
    .a(\D1/n4 [7]),
    .b(\D1/PixelCount [7]),
    .c(\D1/FrameFlag ),
    .d(\D1/mux3_b0_sel_is_0_o ),
    .o(\D1/n8 [7]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u262 (
    .a(\D1/n4 [6]),
    .b(\D1/PixelCount [6]),
    .c(\D1/FrameFlag ),
    .d(\D1/mux3_b0_sel_is_0_o ),
    .o(\D1/n8 [6]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u263 (
    .a(\D1/n4 [5]),
    .b(\D1/PixelCount [5]),
    .c(\D1/FrameFlag ),
    .d(\D1/mux3_b0_sel_is_0_o ),
    .o(\D1/n8 [5]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u264 (
    .a(\D1/n4 [4]),
    .b(\D1/PixelCount [4]),
    .c(\D1/FrameFlag ),
    .d(\D1/mux3_b0_sel_is_0_o ),
    .o(\D1/n8 [4]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u265 (
    .a(\D1/n4 [3]),
    .b(\D1/PixelCount [3]),
    .c(\D1/FrameFlag ),
    .d(\D1/mux3_b0_sel_is_0_o ),
    .o(\D1/n8 [3]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u266 (
    .a(\D1/n4 [2]),
    .b(\D1/PixelCount [2]),
    .c(\D1/FrameFlag ),
    .d(\D1/mux3_b0_sel_is_0_o ),
    .o(\D1/n8 [2]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u267 (
    .a(\D1/n4 [1]),
    .b(\D1/PixelCount [1]),
    .c(\D1/FrameFlag ),
    .d(\D1/mux3_b0_sel_is_0_o ),
    .o(\D1/n8 [1]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u268 (
    .a(\D1/n4 [15]),
    .b(\D1/PixelCount [15]),
    .c(\D1/FrameFlag ),
    .d(\D1/mux3_b0_sel_is_0_o ),
    .o(\D1/n8 [15]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u269 (
    .a(\D1/n4 [14]),
    .b(\D1/PixelCount [14]),
    .c(\D1/FrameFlag ),
    .d(\D1/mux3_b0_sel_is_0_o ),
    .o(\D1/n8 [14]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u270 (
    .a(\D1/n4 [13]),
    .b(\D1/PixelCount [13]),
    .c(\D1/FrameFlag ),
    .d(\D1/mux3_b0_sel_is_0_o ),
    .o(\D1/n8 [13]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u271 (
    .a(\D1/n4 [12]),
    .b(\D1/PixelCount [12]),
    .c(\D1/FrameFlag ),
    .d(\D1/mux3_b0_sel_is_0_o ),
    .o(\D1/n8 [12]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u272 (
    .a(\D1/n4 [11]),
    .b(\D1/PixelCount [11]),
    .c(\D1/FrameFlag ),
    .d(\D1/mux3_b0_sel_is_0_o ),
    .o(\D1/n8 [11]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u273 (
    .a(\D1/n4 [10]),
    .b(\D1/PixelCount [10]),
    .c(\D1/FrameFlag ),
    .d(\D1/mux3_b0_sel_is_0_o ),
    .o(\D1/n8 [10]));
  AL_MAP_LUT4 #(
    .EQN("(D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'hac00))
    _al_u274 (
    .a(\D1/n4 [0]),
    .b(\D1/PixelCount [0]),
    .c(\D1/FrameFlag ),
    .d(\D1/mux3_b0_sel_is_0_o ),
    .o(\D1/n8 [0]));
  AL_MAP_LUT5 #(
    .EQN("~((D*C)*~((B*A))*~(E)+(D*C)*(B*A)*~(E)+~((D*C))*(B*A)*E+(D*C)*(B*A)*E)"),
    .INIT(32'h77770fff))
    _al_u275 (
    .a(\U4/n31 ),
    .b(\U4/n33 ),
    .c(\U4/n37 ),
    .d(\U4/n39 ),
    .e(\U4/AddrCtrl [0]),
    .o(\U4/mux10_b0_sel_is_0_o ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~(B*A))"),
    .INIT(16'h7000))
    _al_u276 (
    .a(\U4/n37 ),
    .b(\U4/n39 ),
    .c(\U4/n23 ),
    .d(\U4/n43 ),
    .o(_al_u276_o));
  AL_MAP_LUT4 #(
    .EQN("~((B*A)*~(C)*~(D)+(B*A)*C*~(D)+~((B*A))*C*D+(B*A)*C*D)"),
    .INIT(16'h0f77))
    _al_u277 (
    .a(\U4/n33 ),
    .b(\U4/n31 ),
    .c(\U4/n27 ),
    .d(\U4/AddrCtrl [0]),
    .o(_al_u277_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*A))"),
    .INIT(8'h0d))
    _al_u278 (
    .a(\U4/n27 ),
    .b(\U4/AddrCtrl [0]),
    .c(\U4/LCD_Ctrl_Reg [4]),
    .o(_al_u278_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~(~B*A))"),
    .INIT(16'hd000))
    _al_u279 (
    .a(\U4/mux10_b0_sel_is_0_o ),
    .b(_al_u276_o),
    .c(_al_u277_o),
    .d(_al_u278_o),
    .o(_al_u279_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u280 (
    .a(i8080_D_pad[7]),
    .b(\U4/LCD_Ctrl_Reg [4]),
    .c(_al_u279_o),
    .o(FIFO_DI[7]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u281 (
    .a(i8080_D_pad[6]),
    .b(\U4/LCD_Ctrl_Reg [4]),
    .c(_al_u279_o),
    .o(FIFO_DI[6]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u282 (
    .a(i8080_D_pad[5]),
    .b(\U4/LCD_Ctrl_Reg [4]),
    .c(_al_u279_o),
    .o(FIFO_DI[5]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~(B*A)))"),
    .INIT(16'h8f00))
    _al_u283 (
    .a(\U4/mux10_b0_sel_is_0_o ),
    .b(_al_u276_o),
    .c(_al_u277_o),
    .d(_al_u278_o),
    .o(_al_u283_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u284 (
    .a(i8080_D_pad[2]),
    .b(\U4/LCD_Ctrl_Reg [4]),
    .c(_al_u283_o),
    .o(FIFO_DI[2]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u285 (
    .a(i8080_D_pad[1]),
    .b(\U4/LCD_Ctrl_Reg [4]),
    .c(_al_u283_o),
    .o(FIFO_DI[1]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u286 (
    .a(i8080_D_pad[0]),
    .b(\U4/LCD_Ctrl_Reg [4]),
    .c(_al_u283_o),
    .o(FIFO_DI[0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*B*~A))"),
    .INIT(16'h00bf))
    _al_u287 (
    .a(\U4/AddrCtrl [0]),
    .b(\U4/n37 ),
    .c(\U4/n39 ),
    .d(_al_u276_o),
    .o(_al_u287_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~(~C*~(~D*~(B*A))))"),
    .INIT(32'hf0f70000))
    _al_u288 (
    .a(\U4/n31 ),
    .b(\U4/n33 ),
    .c(\U4/n27 ),
    .d(_al_u287_o),
    .e(_al_u278_o),
    .o(_al_u288_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u289 (
    .a(\U4/LCD_Ctrl_Reg [4]),
    .b(i8080_D_pad[4]),
    .c(_al_u288_o),
    .o(FIFO_DI[4]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(B*A))"),
    .INIT(8'hf8))
    _al_u290 (
    .a(\U4/LCD_Ctrl_Reg [4]),
    .b(i8080_D_pad[3]),
    .c(_al_u288_o),
    .o(FIFO_DI[3]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u291 (
    .a(FIFO_EMPTY),
    .o(\D1/n28 ));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u292 (
    .a(FIFO_EMPTY),
    .o(LCD_B_pad[2]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u293 (
    .a(\FIFO0/logic_fifo_full ),
    .o(\FIFO0/logic_fifo_full_neg ));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u294 (
    .a(LED_pad[0]),
    .o(\U1/n2 ));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u295 (
    .a(LED_pad[1]),
    .o(\U2/n2 ));
  EF2_PHY_SPAD #(
    //.LOCATION("P54"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u64 (
    .do({open_n511,LCD_B_pad[7]}),
    .ts(1'b1),
    .opad(LCD_B[7]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(21)
  EF2_PHY_SPAD #(
    //.LOCATION("P53"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u65 (
    .do({open_n520,LCD_B_pad[6]}),
    .ts(1'b1),
    .opad(LCD_B[6]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(21)
  EF2_PHY_SPAD #(
    //.LOCATION("P52"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u66 (
    .do({open_n529,LCD_B_pad[5]}),
    .ts(1'b1),
    .opad(LCD_B[5]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(21)
  EF2_PHY_SPAD #(
    //.LOCATION("P51"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u67 (
    .do({open_n538,LCD_B_pad[4]}),
    .ts(1'b1),
    .opad(LCD_B[4]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(21)
  EF2_PHY_PAD #(
    //.LOCATION("P49"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u68 (
    .do({open_n546,open_n547,open_n548,LCD_B_pad[3]}),
    .opad(LCD_B[3]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(21)
  EF2_PHY_PAD #(
    //.LOCATION("P48"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u69 (
    .do({open_n569,open_n570,open_n571,LCD_B_pad[2]}),
    .opad(LCD_B[2]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(21)
  EF2_PHY_PAD #(
    //.LOCATION("P47"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u70 (
    .do({open_n592,open_n593,open_n594,LCD_B_pad[2]}),
    .opad(LCD_B[1]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(21)
  EF2_PHY_PAD #(
    //.LOCATION("P45"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u71 (
    .do({open_n615,open_n616,open_n617,LCD_B_pad[2]}),
    .opad(LCD_B[0]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(21)
  EF2_PHY_SPAD #(
    //.LOCATION("P62"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u72 (
    .do({open_n639,LCD_CLK_pad}),
    .ts(1'b1),
    .opad(LCD_CLK));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(15)
  EF2_PHY_SPAD #(
    //.LOCATION("P60"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u73 (
    .do({open_n648,LCD_DEN_pad}),
    .ts(1'b1),
    .opad(LCD_DEN));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(18)
  EF2_PHY_PAD #(
    //.LOCATION("P43"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u74 (
    .do({open_n656,open_n657,open_n658,LCD_G_pad[7]}),
    .opad(LCD_G[7]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(20)
  EF2_PHY_PAD #(
    //.LOCATION("P42"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u75 (
    .do({open_n679,open_n680,open_n681,LCD_G_pad[6]}),
    .opad(LCD_G[6]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(20)
  EF2_PHY_PAD #(
    //.LOCATION("P41"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u76 (
    .do({open_n702,open_n703,open_n704,LCD_G_pad[5]}),
    .opad(LCD_G[5]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(20)
  EF2_PHY_PAD #(
    //.LOCATION("P40"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u77 (
    .do({open_n725,open_n726,open_n727,LCD_G_pad[4]}),
    .opad(LCD_G[4]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(20)
  EF2_PHY_PAD #(
    //.LOCATION("P39"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u78 (
    .do({open_n748,open_n749,open_n750,LCD_G_pad[3]}),
    .opad(LCD_G[3]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(20)
  EF2_PHY_PAD #(
    //.LOCATION("P38"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u79 (
    .do({open_n771,open_n772,open_n773,LCD_G_pad[2]}),
    .opad(LCD_G[2]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(20)
  EF2_PHY_PAD #(
    //.LOCATION("P37"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u80 (
    .do({open_n794,open_n795,open_n796,LCD_B_pad[2]}),
    .opad(LCD_G[1]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(20)
  EF2_PHY_PAD #(
    //.LOCATION("P36"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u81 (
    .do({open_n817,open_n818,open_n819,LCD_B_pad[2]}),
    .opad(LCD_G[0]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(20)
  EF2_PHY_SPAD #(
    //.LOCATION("P58"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u82 (
    .do({open_n841,LCD_HYNC_pad}),
    .ts(1'b1),
    .opad(LCD_HYNC));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(16)
  EF2_PHY_PAD #(
    //.LOCATION("P35"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u83 (
    .do({open_n849,open_n850,open_n851,LCD_R_pad[7]}),
    .opad(LCD_R[7]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(19)
  EF2_PHY_PAD #(
    //.LOCATION("P34"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u84 (
    .do({open_n872,open_n873,open_n874,LCD_R_pad[6]}),
    .opad(LCD_R[6]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(19)
  EF2_PHY_PAD #(
    //.LOCATION("P32"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u85 (
    .do({open_n895,open_n896,open_n897,LCD_R_pad[5]}),
    .opad(LCD_R[5]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(19)
  EF2_PHY_PAD #(
    //.LOCATION("P31"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u86 (
    .do({open_n918,open_n919,open_n920,LCD_R_pad[4]}),
    .opad(LCD_R[4]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(19)
  EF2_PHY_PAD #(
    //.LOCATION("P30"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u87 (
    .do({open_n941,open_n942,open_n943,LCD_R_pad[3]}),
    .opad(LCD_R[3]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(19)
  EF2_PHY_PAD #(
    //.LOCATION("P29"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u88 (
    .do({open_n964,open_n965,open_n966,1'b1}),
    .opad(LCD_R[2]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(19)
  EF2_PHY_PAD #(
    //.LOCATION("P28"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u89 (
    .do({open_n987,open_n988,open_n989,1'b1}),
    .opad(LCD_R[1]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(19)
  EF2_PHY_PAD #(
    //.LOCATION("P27"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u90 (
    .do({open_n1010,open_n1011,open_n1012,1'b1}),
    .opad(LCD_R[0]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(19)
  EF2_PHY_SPAD #(
    //.LOCATION("P59"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u91 (
    .do({open_n1034,LCD_SYNC_pad}),
    .ts(1'b1),
    .opad(LCD_SYNC));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(17)
  EF2_PHY_SPAD #(
    //.LOCATION("P63"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u92 (
    .do({open_n1043,LED_pad[1]}),
    .ts(1'b1),
    .opad(LED[1]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(6)
  EF2_PHY_SPAD #(
    //.LOCATION("P64"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u93 (
    .do({open_n1052,LED_pad[0]}),
    .ts(1'b1),
    .opad(LED[0]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(6)
  EF2_PHY_SPAD #(
    //.LOCATION("P4"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u94 (
    .ipad(clk),
    .ts(1'b1),
    .di(clk_pad));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(3)
  EF2_PHY_SPAD #(
    //.LOCATION("P10"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS18"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u95 (
    .ipad(i8080_CS),
    .ts(1'b1),
    .di(i8080_CS_pad));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("P16"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS18"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u96 (
    .ipad(i8080_D[7]),
    .ts(1'b1),
    .di(i8080_D_pad[7]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(12)
  EF2_PHY_SPAD #(
    //.LOCATION("P17"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS18"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u97 (
    .ipad(i8080_D[6]),
    .ts(1'b1),
    .di(i8080_D_pad[6]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(12)
  EF2_PHY_SPAD #(
    //.LOCATION("P18"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS18"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u98 (
    .ipad(i8080_D[5]),
    .ts(1'b1),
    .di(i8080_D_pad[5]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(12)
  EF2_PHY_SPAD #(
    //.LOCATION("P21"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS18"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u99 (
    .ipad(i8080_D[2]),
    .ts(1'b1),
    .di(i8080_D_pad[2]));  // E:/Fpga_Prj/Anlogic/LCD_8080ToRGB/source/TOP.v(12)
  EF2_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();

endmodule 

module reg_ar_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(enout),
    .reset(reset),
    .set(set),
    .q(q));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

